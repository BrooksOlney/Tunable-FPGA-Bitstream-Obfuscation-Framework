module ks_apex4_qmap_map (sk, i_0_, i_1_, i_2_, i_6_, i_7_, i_8_, i_3_, i_4_, i_5_, o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_);

	input i_0_;
	input i_1_;
	input i_2_;
	input i_6_;
	input i_7_;
	input i_8_;
	input i_3_;
	input i_4_;
	input i_5_;
	output o_0_;
	output o_1_;
	output o_2_;
	output o_3_;
	output o_4_;
	output o_5_;
	output o_6_;
	output o_7_;
	output o_8_;
	output o_9_;
	output o_10_;
	output o_11_;
	output o_12_;
	output o_13_;
	output o_14_;
	output o_15_;
	output o_16_;
	output o_17_;
	output o_18_;

	input [127 : 0] sk /* synthesis noprune */;


	wire gnd, g82, g199, g263, g320, g356, g395, g418, g437, g454, g467, g490, g510, g520, g523, g532, g537, g540, g542, g1, g2;
	wire g3, g4, g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g20, g21, g22, g23;
	wire g24, g25, g26, g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37, g38, g39, g40, g41, g42, g43, g44;
	wire g45, g46, g47, g48, g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59, g60, g61, g62, g63, g64, g65;
	wire g66, g67, g68, g69, g70, g71, g72, g73, g74, g75, g76, g77, g78, g79, g80, g81, g83, g84, g85, g86, g87;
	wire g88, g89, g90, g91, g92, g93, g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104, g105, g106, g107, g108;
	wire g109, g110, g111, g112, g113, g114, g115, g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126, g127, g128, g129;
	wire g130, g131, g683, g132, g694, g133, g134, g135, g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146, g147, g148;
	wire g149, g150, g151, g152, g670, g153, g154, g155, g156, g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167, g168;
	wire g169, g170, g171, g172, g173, g174, g175, g176, g177, g178, g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189;
	wire g190, g657, g191, g192, g193, g194, g195, g196, g197, g198, g200, g201, g202, g203, g204, g205, g206, g207, g208, g209, g644;
	wire g210, g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221, g222, g223, g224, g225, g226, g227, g228, g229, g230;
	wire g231, g232, g631, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242, g243, g244, g245, g246, g247, g248, g249, g250;
	wire g251, g252, g253, g254, g255, g256, g257, g258, g259, g260, g261, g262, g264, g265, g266, g267, g268, g269, g270, g271, g272;
	wire g273, g274, g275, g276, g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287, g288, g289, g290, g291, g292, g293;
	wire g294, g295, g296, g297, g298, g299, g300, g301, g302, g303, g304, g305, g607, g306, g307, g308, g309, g310, g311, g312, g313;
	wire g314, g315, g316, g317, g318, g319, g618, g321, g322, g596, g323, g324, g325, g326, g327, g328, g329, g330, g331, g332, g333;
	wire g334, g335, g336, g337, g338, g339, g340, g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351, g352, g353, g354;
	wire g355, g357, g358, g359, g360, g361, g362, g363, g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374, g375, g376;
	wire g377, g378, g379, g380, g381, g382, g383, g384, g385, g386, g387, g388, g389, g390, g391, g392, g583, g393, g394, g396, g397;
	wire g398, g399, g400, g401, g402, g403, g404, g405, g406, g407, g408, g409, g410, g411, g412, g413, g414, g415, g416, g417, g419;
	wire g420, g421, g422, g572, g423, g424, g425, g426, g427, g428, g429, g430, g431, g432, g433, g434, g435, g436, g438, g439, g440;
	wire g441, g442, g443, g444, g445, g446, g447, g448, g449, g559, g450, g451, g452, g453, g455, g456, g457, g458, g459, g460, g461;
	wire g462, g463, g464, g465, g466, g468, g469, g470, g471, g472, g473, g474, g475, g476, g477, g478, g549, g479, g480, g481, g482;
	wire g483, g484, g485, g486, g487, g488, g489, g491, g492, g493, g494, g495, g496, g497, g498, g499, g500, g501, g502, g503, g504;
	wire g505, g506, g507, g508, g509, g511, g512, g513, g514, g515, g516, g517, g543, g518, g519, g521, g522, g524, g525, g526, g527;
	wire g528, g529, g530, g531, g533, g534, g535, g536, g538, g539, g541, g544, g545, g546, g547, g548, g550, g551, g552, g554, g553;
	wire g555, g556, g557, g558, g560, g561, g562, g565, g563, g564, g568, g569, g566, g567, g570, g571, g573, g574, g575, g578, g576;
	wire g577, g580, g581, g579, g582, g584, g585, g586, g589, g587, g588, g592, g593, g590, g591, g594, g595, g597, g598, g599, g601;
	wire g600, g604, g602, g603, g605, g606, g608, g609, g610, g612, g611, g615, g613, g614, g616, g617, g619, g620, g621, g624, g622;
	wire g623, g627, g628, g625, g626, g629, g630, g632, g633, g634, g637, g635, g636, g640, g641, g638, g639, g642, g643, g645, g646;
	wire g647, g650, g648, g649, g653, g654, g651, g652, g655, g656, g658, g659, g660, g663, g661, g662, g666, g667, g664, g665, g668;
	wire g669, g671, g672, g673, g676, g674, g675, g679, g680, g677, g678, g681, g682, g684, g685, g686, g689, g687, g688, g691, g692;
	wire g690, g693, g695, g696, g697, g699, g698, g702, g700, g701, g703, g704;

	assign o_0_ = (((sk[0]) & (gnd)));
	assign o_1_ = (((sk[1]) & (!g82)));
	assign o_2_ = (((sk[2]) & (!g199)));
	assign o_3_ = (((sk[3]) & (!g263)));
	assign o_4_ = (((sk[4]) & (!g320)));
	assign o_5_ = (((sk[5]) & (!g356)));
	assign o_6_ = (((sk[6]) & (!g395)));
	assign o_7_ = (((sk[7]) & (!g418)));
	assign o_8_ = (((sk[8]) & (!g437)));
	assign o_9_ = (((sk[9]) & (!g454)));
	assign o_10_ = (((sk[10]) & (!g467)));
	assign o_11_ = (((sk[11]) & (!g490)));
	assign o_12_ = (((sk[12]) & (!g510)));
	assign o_13_ = (((sk[13]) & (!g520)));
	assign o_14_ = (((sk[14]) & (!g523)));
	assign o_15_ = (((sk[15]) & (!g532)));
	assign o_16_ = (((sk[16]) & (!g537)));
	assign o_17_ = (((sk[17]) & (!g540)));
	assign o_18_ = (((sk[18]) & (!g542)));
	assign g1 = (((!i_0_) & (sk[19]) & (!i_1_) & (!i_2_)) + ((i_0_) & (!sk[19]) & (i_1_) & (!i_2_)) + ((!i_0_) & (sk[19]) & (!i_1_) & (i_2_)));
	assign g2 = (((i_6_) & (i_7_) & (!sk[20]) & (!i_8_)) + ((i_6_) & (!i_7_) & (sk[20]) & (!i_8_)));
	assign g3 = (((i_3_) & (!sk[21]) & (i_4_) & (!i_5_)) + ((!i_3_) & (sk[21]) & (i_4_) & (!i_5_)));
	assign g4 = (((g2) & (!sk[22]) & (g3)));
	assign g5 = (((!i_3_) & (sk[23]) & (i_4_)) + ((i_3_) & (!sk[23]) & (i_4_)));
	assign g6 = (((i_6_) & (!sk[24]) & (i_7_) & (!i_8_)) + ((i_6_) & (sk[24]) & (!i_7_) & (i_8_)));
	assign g7 = (((!sk[25]) & (g1) & (g6)) + ((sk[25]) & (!g1) & (g6)));
	assign g8 = (((i_6_) & (i_7_) & (!sk[26]) & (!i_8_)) + ((!i_6_) & (i_7_) & (sk[26]) & (i_8_)));
	assign g9 = (((!sk[27]) & (g8) & (g1)) + ((sk[27]) & (g8) & (!g1)));
	assign g10 = (((i_5_) & (g5) & (!sk[28]) & (!g7) & (!g9)) + ((i_5_) & (g5) & (!sk[28]) & (g7) & (!g9)) + ((!i_5_) & (g5) & (sk[28]) & (!g7) & (g9)));
	assign g11 = (((!sk[29]) & (!i_3_) & (!i_4_) & (i_5_)) + ((sk[29]) & (!i_3_) & (!i_4_) & (!i_5_)) + ((!sk[29]) & (i_3_) & (!i_4_) & (i_5_)) + ((!sk[29]) & (!i_3_) & (i_4_) & (i_5_)));
	assign g12 = (((!i_6_) & (!sk[30]) & (!i_7_) & (i_8_)) + ((!i_6_) & (sk[30]) & (i_7_) & (!i_8_)));
	assign g13 = (((!i_0_) & (!sk[31]) & (!i_1_) & (i_2_)) + ((!i_0_) & (sk[31]) & (!i_1_) & (!i_2_)) + ((!i_0_) & (sk[31]) & (!i_1_) & (!i_2_)));
	assign g14 = (((i_7_) & (!sk[32]) & (i_8_)) + ((!i_7_) & (!sk[32]) & (i_8_)));
	assign g15 = (((!i_4_) & (!sk[33]) & (!i_5_) & (i_6_)) + ((i_4_) & (sk[33]) & (i_5_) & (!i_6_)));
	assign g16 = (((!sk[34]) & (!g14) & (g15)) + ((!sk[34]) & (g14) & (g15)));
	assign g17 = (((!sk[35]) & (!i_3_) & (!i_0_) & (i_2_)) + ((sk[35]) & (i_3_) & (i_0_) & (!i_2_)));
	assign g18 = (((!sk[36]) & (!g16) & (g17)) + ((!sk[36]) & (g16) & (g17)));
	assign g19 = (((!sk[37]) & (!g11) & (g12) & (!g13) & (!g18)) + ((!sk[37]) & (!g11) & (!g12) & (g13) & (!g18)) + ((!sk[37]) & (!g11) & (!g12) & (g13) & (!g18)) + ((sk[37]) & (!g11) & (!g12) & (!g13) & (!g18)) + ((!sk[37]) & (g11) & (g12) & (!g13) & (!g18)));
	assign g20 = (((!g1) & (!sk[38]) & (g4) & (!g10) & (!g19)) + ((!g1) & (!sk[38]) & (!g4) & (g10) & (!g19)) + ((!g1) & (sk[38]) & (!g4) & (!g10) & (g19)) + ((g1) & (!sk[38]) & (g4) & (!g10) & (g19)));
	assign g21 = (((!i_3_) & (!sk[39]) & (!i_4_) & (i_5_)) + ((!i_3_) & (sk[39]) & (!i_4_) & (!i_5_)) + ((!i_3_) & (!sk[39]) & (!i_4_) & (i_5_)) + ((!i_3_) & (!sk[39]) & (i_4_) & (i_5_)));
	assign g22 = (((!g21) & (!sk[40]) & (g2)) + ((!g21) & (!sk[40]) & (g2)));
	assign g23 = (((!i_6_) & (!i_7_) & (!sk[41]) & (i_8_)) + ((!i_6_) & (!i_7_) & (sk[41]) & (!i_8_)) + ((!i_6_) & (!i_7_) & (sk[41]) & (!i_8_)));
	assign g24 = (((!i_0_) & (!sk[42]) & (!i_1_) & (i_2_)) + ((!i_0_) & (sk[42]) & (!i_1_) & (!i_2_)) + ((i_0_) & (!sk[42]) & (!i_1_) & (i_2_)) + ((!i_0_) & (!sk[42]) & (!i_1_) & (i_2_)));
	assign g25 = (((!i_0_) & (!i_1_) & (!sk[43]) & (i_2_)) + ((i_0_) & (!i_1_) & (sk[43]) & (!i_2_)) + ((!i_0_) & (!i_1_) & (sk[43]) & (!i_2_)));
	assign g26 = (((!g11) & (!sk[44]) & (g25)) + ((!g11) & (sk[44]) & (!g25)));
	assign g27 = (((!i_0_) & (!sk[45]) & (!i_1_) & (i_2_)) + ((!i_0_) & (sk[45]) & (!i_1_) & (!i_2_)) + ((!i_0_) & (!sk[45]) & (!i_1_) & (i_2_)) + ((!i_0_) & (!sk[45]) & (!i_1_) & (i_2_)));
	assign g28 = (((!sk[46]) & (!i_6_) & (!i_7_) & (i_8_)) + ((!sk[46]) & (i_6_) & (i_7_) & (i_8_)));
	assign g29 = (((!g28) & (!sk[47]) & (g1)) + ((g28) & (sk[47]) & (!g1)));
	assign g30 = (((g11) & (!g27) & (!g21) & (!g6) & (!sk[48]) & (!g29)) + ((!g11) & (!g27) & (g21) & (!g6) & (!sk[48]) & (!g29)) + ((!g11) & (g27) & (!g21) & (g6) & (!sk[48]) & (!g29)) + ((!g11) & (!g27) & (!g21) & (!g6) & (sk[48]) & (g29)) + ((!g11) & (!g27) & (!g21) & (g6) & (sk[48]) & (!g29)));
	assign g31 = (((g22) & (!g23) & (!sk[49]) & (!g24) & (!g26) & (!g30)) + ((!g22) & (!g23) & (!sk[49]) & (g24) & (!g26) & (!g30)) + ((!g22) & (g23) & (!sk[49]) & (!g24) & (g26) & (!g30)) + ((!g22) & (g23) & (!sk[49]) & (g24) & (!g26) & (!g30)) + ((!g22) & (!g23) & (!sk[49]) & (g24) & (!g26) & (!g30)) + ((!g22) & (!g23) & (sk[49]) & (!g24) & (!g26) & (!g30)) + ((!g22) & (g23) & (!sk[49]) & (!g24) & (g26) & (!g30)));
	assign g32 = (((!i_3_) & (!sk[50]) & (!i_4_) & (i_5_)) + ((!i_3_) & (sk[50]) & (!i_4_) & (!i_5_)));
	assign g33 = (((!sk[51]) & (!g24) & (g3)) + ((!sk[51]) & (!g24) & (g3)));
	assign g34 = (((!g11) & (!g27) & (!g6) & (!g23) & (!g32) & (g33)) + ((!g11) & (!g27) & (!g6) & (!g23) & (!g32) & (!g33)) + ((!g11) & (!g27) & (g6) & (!g23) & (g32) & (!g33)));
	assign g35 = (((!i_6_) & (!sk[53]) & (!i_7_) & (i_8_)) + ((!i_6_) & (sk[53]) & (!i_7_) & (!i_8_)));
	assign g36 = (((!i_3_) & (!sk[54]) & (!i_4_) & (i_5_)) + ((!i_3_) & (sk[54]) & (!i_4_) & (!i_5_)) + ((!i_3_) & (sk[54]) & (i_4_) & (!i_5_)));
	assign g37 = (((!sk[55]) & (!i_6_) & (i_7_)) + ((sk[55]) & (!i_6_) & (!i_7_)));
	assign g38 = (((!i_3_) & (!sk[56]) & (!i_4_) & (i_5_)) + ((!i_3_) & (sk[56]) & (!i_4_) & (!i_5_)) + ((i_3_) & (!sk[56]) & (!i_4_) & (i_5_)) + ((!i_3_) & (!sk[56]) & (!i_4_) & (i_5_)));
	assign g39 = (((g11) & (!sk[57]) & (!g27) & (!g2) & (!g37) & (!g38)) + ((!g11) & (!sk[57]) & (!g27) & (g2) & (!g37) & (!g38)) + ((!g11) & (!sk[57]) & (!g27) & (g2) & (!g37) & (!g38)) + ((!g11) & (!sk[57]) & (g27) & (!g2) & (g37) & (!g38)) + ((!g11) & (sk[57]) & (!g27) & (!g2) & (g37) & (!g38)));
	assign g40 = (((!g35) & (!sk[58]) & (g1) & (!g36) & (!g39)) + ((!g35) & (!sk[58]) & (!g1) & (g36) & (!g39)) + ((!g35) & (!sk[58]) & (g1) & (!g36) & (!g39)) + ((!g35) & (!sk[58]) & (!g1) & (g36) & (!g39)) + ((!g35) & (sk[58]) & (!g1) & (!g36) & (!g39)));
	assign g41 = (((!g27) & (!sk[59]) & (g35)) + ((!g27) & (!sk[59]) & (g35)));
	assign g42 = (((!i_0_) & (!i_1_) & (!sk[60]) & (i_2_)) + ((i_0_) & (!i_1_) & (!sk[60]) & (i_2_)));
	assign g43 = (((!sk[61]) & (!g21) & (!g28) & (g42)) + ((!sk[61]) & (!g21) & (g28) & (g42)));
	assign g44 = (((!g11) & (!sk[62]) & (g41) & (!g43) & (!g3)) + ((!g11) & (!sk[62]) & (!g41) & (g43) & (!g3)) + ((!g11) & (sk[62]) & (!g41) & (!g43) & (!g3)) + ((g11) & (!sk[62]) & (g41) & (!g43) & (!g3)));
	assign g45 = (((!sk[63]) & (!i_3_) & (!i_4_) & (i_5_)) + ((sk[63]) & (!i_3_) & (!i_4_) & (!i_5_)) + ((sk[63]) & (!i_3_) & (!i_4_) & (!i_5_)));
	assign g46 = (((!sk[64]) & (!g25) & (g45)) + ((sk[64]) & (!g25) & (!g45)));
	assign g47 = (((!i_7_) & (!sk[65]) & (i_8_)) + ((!i_7_) & (!sk[65]) & (i_8_)));
	assign g48 = (((!sk[66]) & (!i_6_) & (g47)) + ((!sk[66]) & (!i_6_) & (g47)));
	assign g49 = (((!g32) & (!sk[67]) & (g13)) + ((g32) & (sk[67]) & (!g13)));
	assign g50 = (((!i_4_) & (!sk[68]) & (i_5_)) + ((!i_4_) & (!sk[68]) & (i_5_)));
	assign g51 = (((!i_3_) & (!i_0_) & (!sk[69]) & (i_2_)) + ((!i_3_) & (i_0_) & (sk[69]) & (!i_2_)));
	assign g52 = (((!sk[70]) & (!g50) & (g51)) + ((!sk[70]) & (g50) & (g51)));
	assign g53 = (((!sk[71]) & (g8) & (!g46) & (!g48) & (!g49) & (!g52)) + ((!sk[71]) & (!g8) & (!g46) & (g48) & (!g49) & (!g52)) + ((sk[71]) & (!g8) & (!g46) & (!g48) & (!g49) & (!g52)) + ((!sk[71]) & (g8) & (!g46) & (!g48) & (!g49) & (!g52)) + ((!sk[71]) & (!g8) & (g46) & (!g48) & (g49) & (!g52)) + ((!sk[71]) & (!g8) & (!g46) & (g48) & (!g49) & (!g52)) + ((!sk[71]) & (!g8) & (!g46) & (g48) & (!g49) & (!g52)));
	assign g54 = (((i_4_) & (!sk[72]) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_8_)) + ((!i_4_) & (!sk[72]) & (!i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((!i_4_) & (!sk[72]) & (i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((i_4_) & (!sk[72]) & (!i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((!i_4_) & (sk[72]) & (!i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((!i_4_) & (!sk[72]) & (i_5_) & (i_6_) & (i_7_) & (!i_8_)));
	assign g55 = (((!sk[73]) & (g50) & (!g42) & (!g1) & (!g12) & (!g22)) + ((!sk[73]) & (!g50) & (!g42) & (g1) & (!g12) & (!g22)) + ((!sk[73]) & (!g50) & (g42) & (!g1) & (g12) & (!g22)) + ((!sk[73]) & (g50) & (!g42) & (!g1) & (g12) & (!g22)) + ((sk[73]) & (!g50) & (g42) & (!g1) & (!g12) & (g22)));
	assign g56 = (((!i_3_) & (!sk[74]) & (g1) & (!g54) & (!g55)) + ((!i_3_) & (!sk[74]) & (!g1) & (g54) & (!g55)) + ((!i_3_) & (!sk[74]) & (g1) & (!g54) & (!g55)) + ((!i_3_) & (sk[74]) & (!g1) & (!g54) & (!g55)) + ((!i_3_) & (!sk[74]) & (!g1) & (g54) & (!g55)));
	assign g57 = (((!i_3_) & (!i_1_) & (!sk[75]) & (i_2_)) + ((i_3_) & (!i_1_) & (!sk[75]) & (i_2_)));
	assign g58 = (((!sk[76]) & (!i_4_) & (i_5_) & (!g57) & (!g6)) + ((!sk[76]) & (!i_4_) & (!i_5_) & (g57) & (!g6)) + ((!sk[76]) & (i_4_) & (i_5_) & (g57) & (g6)));
	assign g59 = (((!i_3_) & (!i_4_) & (!sk[77]) & (i_5_)) + ((!i_3_) & (!i_4_) & (sk[77]) & (!i_5_)) + ((!i_3_) & (!i_4_) & (!sk[77]) & (i_5_)) + ((!i_3_) & (!i_4_) & (!sk[77]) & (i_5_)));
	assign g60 = (((!sk[78]) & (!i_6_) & (i_7_)) + ((!sk[78]) & (i_6_) & (i_7_)));
	assign g61 = (((g42) & (!g58) & (!sk[79]) & (!g59) & (!g13) & (!g60)) + ((!g42) & (!g58) & (!sk[79]) & (g59) & (!g13) & (!g60)) + ((!g42) & (!g58) & (!sk[79]) & (g59) & (!g13) & (!g60)) + ((!g42) & (g58) & (!sk[79]) & (!g59) & (g13) & (!g60)) + ((!g42) & (!g58) & (sk[79]) & (!g59) & (!g13) & (!g60)) + ((!g42) & (!g58) & (sk[79]) & (!g59) & (g13) & (!g60)));
	assign g62 = (((!sk[80]) & (g40) & (!g44) & (!g53) & (!g56) & (!g61)) + ((!sk[80]) & (!g40) & (!g44) & (g53) & (!g56) & (!g61)) + ((!sk[80]) & (!g40) & (g44) & (!g53) & (g56) & (!g61)) + ((!sk[80]) & (g40) & (g44) & (g53) & (g56) & (g61)));
	assign g63 = (((!i_7_) & (!sk[81]) & (i_8_)) + ((!i_7_) & (sk[81]) & (!i_8_)));
	assign g64 = (((!i_4_) & (!sk[82]) & (!i_5_) & (i_6_)) + ((i_4_) & (sk[82]) & (!i_5_) & (!i_6_)));
	assign g65 = (((!i_3_) & (!sk[83]) & (i_0_) & (!i_1_) & (!g64)) + ((!i_3_) & (!sk[83]) & (!i_0_) & (i_1_) & (!g64)) + ((i_3_) & (!sk[83]) & (i_0_) & (!i_1_) & (g64)));
	assign g66 = (((!sk[84]) & (g42) & (!g45) & (!g23) & (!g36) & (!g29)) + ((!sk[84]) & (!g42) & (!g45) & (g23) & (!g36) & (!g29)) + ((!sk[84]) & (g42) & (!g45) & (!g23) & (!g36) & (!g29)) + ((!sk[84]) & (!g42) & (g45) & (!g23) & (g36) & (!g29)) + ((sk[84]) & (!g42) & (!g45) & (!g23) & (!g36) & (g29)));
	assign g67 = (((!g27) & (!sk[85]) & (g2)) + ((!g27) & (!sk[85]) & (g2)));
	assign g68 = (((g1) & (!sk[86]) & (!g23) & (!g32) & (!g36) & (!g67)) + ((!g1) & (!sk[86]) & (!g23) & (g32) & (!g36) & (!g67)) + ((!g1) & (!sk[86]) & (!g23) & (g32) & (!g36) & (g67)) + ((!g1) & (!sk[86]) & (g23) & (!g32) & (g36) & (!g67)) + ((!g1) & (sk[86]) & (!g23) & (!g32) & (!g36) & (!g67)));
	assign g69 = (((!g42) & (g45) & (!g6) & (!sk[87]) & (!g68)) + ((!g42) & (!g45) & (g6) & (!sk[87]) & (!g68)) + ((!g42) & (g45) & (!g6) & (!sk[87]) & (!g68)) + ((!g42) & (!g45) & (!g6) & (sk[87]) & (!g68)) + ((!g42) & (!g45) & (!g6) & (sk[87]) & (!g68)));
	assign g70 = (((!g25) & (!sk[88]) & (g32)) + ((!g25) & (!sk[88]) & (g32)));
	assign g71 = (((!g42) & (!sk[89]) & (g59)) + ((g42) & (sk[89]) & (!g59)));
	assign g72 = (((g27) & (!g28) & (!g32) & (!g37) & (!sk[90]) & (!g71)) + ((!g27) & (!g28) & (g32) & (!g37) & (!sk[90]) & (!g71)) + ((!g27) & (g28) & (g32) & (!g37) & (!sk[90]) & (!g71)) + ((!g27) & (g28) & (!g32) & (g37) & (!sk[90]) & (!g71)) + ((!g27) & (!g28) & (!g32) & (g37) & (sk[90]) & (g71)));
	assign g73 = (((!g11) & (!sk[91]) & (g24)) + ((!g11) & (sk[91]) & (!g24)));
	assign g74 = (((!g6) & (!g24) & (!sk[92]) & (g32)) + ((g6) & (!g24) & (!sk[92]) & (g32)));
	assign g75 = (((!g24) & (!sk[93]) & (g59)) + ((!g24) & (sk[93]) & (!g59)));
	assign g76 = (((!g23) & (!sk[94]) & (g73) & (!g74) & (!g75)) + ((!g23) & (!sk[94]) & (!g73) & (g74) & (!g75)) + ((g23) & (sk[94]) & (!g73) & (!g74) & (!g75)) + ((!g23) & (sk[94]) & (!g73) & (!g74) & (!g75)));
	assign g77 = (((!sk[95]) & (!g25) & (g59)) + ((sk[95]) & (!g25) & (!g59)));
	assign g78 = (((!g28) & (!sk[96]) & (g2) & (!g77) & (!g33)) + ((!g28) & (!sk[96]) & (!g2) & (g77) & (!g33)) + ((!g28) & (!sk[96]) & (g2) & (g77) & (!g33)) + ((g28) & (sk[96]) & (!g2) & (!g77) & (g33)));
	assign g79 = (((g6) & (!g70) & (!sk[97]) & (!g72) & (!g76) & (!g78)) + ((!g6) & (!g70) & (!sk[97]) & (g72) & (!g76) & (!g78)) + ((!g6) & (g70) & (!sk[97]) & (!g72) & (g76) & (!g78)) + ((!g6) & (!g70) & (sk[97]) & (!g72) & (g76) & (!g78)) + ((!g6) & (!g70) & (sk[97]) & (!g72) & (g76) & (!g78)));
	assign g80 = (((g21) & (!g8) & (!sk[98]) & (!g24) & (!g69) & (!g79)) + ((!g21) & (!g8) & (!sk[98]) & (g24) & (!g69) & (!g79)) + ((!g21) & (g8) & (!sk[98]) & (!g24) & (g69) & (!g79)) + ((g21) & (!g8) & (!sk[98]) & (!g24) & (g69) & (g79)) + ((!g21) & (!g8) & (!sk[98]) & (g24) & (g69) & (g79)) + ((!g21) & (!g8) & (sk[98]) & (!g24) & (g69) & (g79)));
	assign g81 = (((!g63) & (g65) & (!g66) & (!sk[99]) & (!g80)) + ((!g63) & (!g65) & (g66) & (!sk[99]) & (!g80)) + ((!g63) & (!g65) & (!g66) & (sk[99]) & (g80)) + ((!g63) & (!g65) & (!g66) & (sk[99]) & (g80)));
	assign g82 = (((g20) & (!g31) & (!g34) & (!g62) & (!sk[100]) & (!g81)) + ((!g20) & (!g31) & (g34) & (!g62) & (!sk[100]) & (!g81)) + ((!g20) & (g31) & (!g34) & (g62) & (!sk[100]) & (!g81)) + ((g20) & (g31) & (!g34) & (g62) & (!sk[100]) & (g81)));
	assign g83 = (((g21) & (!g8) & (!sk[101]) & (!g24) & (!g77) & (!g37)) + ((!g21) & (!g8) & (!sk[101]) & (g24) & (!g77) & (!g37)) + ((!g21) & (g8) & (!sk[101]) & (!g24) & (g77) & (!g37)) + ((!g21) & (!g8) & (sk[101]) & (!g24) & (!g77) & (g37)));
	assign g84 = (((!g1) & (!sk[102]) & (g38)) + ((!g1) & (sk[102]) & (!g38)));
	assign g85 = (((!i_4_) & (!i_5_) & (!sk[103]) & (i_6_)) + ((!i_4_) & (!i_5_) & (!sk[103]) & (i_6_)));
	assign g86 = (((!i_3_) & (!i_0_) & (!sk[104]) & (i_2_)) + ((i_3_) & (i_0_) & (!sk[104]) & (i_2_)));
	assign g87 = (((g63) & (!g8) & (!sk[105]) & (!g84) & (!g85) & (!g86)) + ((!g63) & (g8) & (!sk[105]) & (g84) & (!g85) & (!g86)) + ((!g63) & (!g8) & (!sk[105]) & (g84) & (!g85) & (!g86)) + ((!g63) & (g8) & (!sk[105]) & (!g84) & (g85) & (!g86)) + ((g63) & (!g8) & (!sk[105]) & (!g84) & (g85) & (g86)));
	assign g88 = (((!sk[106]) & (!g42) & (g36)) + ((sk[106]) & (g42) & (!g36)));
	assign g89 = (((!sk[107]) & (!g23) & (g3) & (!g29) & (!g88)) + ((!sk[107]) & (!g23) & (!g3) & (g29) & (!g88)) + ((!sk[107]) & (!g23) & (g3) & (g29) & (!g88)) + ((sk[107]) & (!g23) & (!g3) & (!g29) & (g88)));
	assign g90 = (((!g45) & (!sk[108]) & (g6) & (!g13) & (!g89)) + ((!g45) & (!sk[108]) & (!g6) & (g13) & (!g89)) + ((!g45) & (!sk[108]) & (!g6) & (g13) & (!g89)) + ((!g45) & (sk[108]) & (!g6) & (!g13) & (!g89)) + ((g45) & (!sk[108]) & (g6) & (!g13) & (!g89)));
	assign g91 = (((!g36) & (!sk[109]) & (g13)) + ((!g36) & (sk[109]) & (!g13)));
	assign g92 = (((!sk[110]) & (!g42) & (!g12) & (g3)) + ((!sk[110]) & (g42) & (g12) & (g3)));
	assign g93 = (((g41) & (!g45) & (!g48) & (!sk[111]) & (!g91) & (!g92)) + ((!g41) & (!g45) & (g48) & (!sk[111]) & (!g91) & (!g92)) + ((!g41) & (g45) & (!g48) & (!sk[111]) & (g91) & (!g92)) + ((!g41) & (!g45) & (!g48) & (sk[111]) & (!g91) & (!g92)) + ((!g41) & (g45) & (!g48) & (sk[111]) & (!g91) & (!g92)) + ((!g41) & (!g45) & (!g48) & (sk[111]) & (!g91) & (!g92)) + ((!g41) & (g45) & (!g48) & (sk[111]) & (!g91) & (!g92)));
	assign g94 = (((!sk[112]) & (!i_3_) & (!i_0_) & (i_1_)) + ((sk[112]) & (!i_3_) & (i_0_) & (!i_1_)));
	assign g95 = (((g47) & (!sk[113]) & (g94)) + ((!g47) & (!sk[113]) & (g94)));
	assign g96 = (((g85) & (!sk[114]) & (g95)) + ((!g85) & (!sk[114]) & (g95)));
	assign g97 = (((!sk[115]) & (!g27) & (!g23) & (g32)) + ((!sk[115]) & (!g27) & (!g23) & (g32)));
	assign g98 = (((!g24) & (!sk[116]) & (g36)) + ((!g24) & (sk[116]) & (!g36)));
	assign g99 = (((!sk[117]) & (!g25) & (g3)) + ((!sk[117]) & (!g25) & (g3)));
	assign g100 = (((!sk[118]) & (!g3) & (g13)) + ((sk[118]) & (g3) & (!g13)));
	assign g101 = (((!i_6_) & (i_7_) & (!i_8_) & (g98) & (!g99) & (!g100)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g98) & (!g99) & (g100)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g98) & (g99) & (!g100)));
	assign g102 = (((!g8) & (g12) & (!sk[120]) & (!g75) & (!g49)) + ((g8) & (!g12) & (!sk[120]) & (g75) & (!g49)) + ((!g8) & (!g12) & (!sk[120]) & (g75) & (!g49)) + ((!g8) & (g12) & (!sk[120]) & (!g75) & (g49)));
	assign g103 = (((!g28) & (!sk[121]) & (g42) & (!g45) & (!g24)) + ((!g28) & (!sk[121]) & (!g42) & (g45) & (!g24)) + ((g28) & (!sk[121]) & (g42) & (!g45) & (!g24)) + ((g28) & (sk[121]) & (!g42) & (!g45) & (!g24)));
	assign g104 = (((!sk[122]) & (!g21) & (g25) & (!g12) & (!g103)) + ((!sk[122]) & (!g21) & (!g25) & (g12) & (!g103)) + ((!sk[122]) & (!g21) & (g25) & (!g12) & (!g103)) + ((sk[122]) & (!g21) & (!g25) & (!g12) & (!g103)) + ((!sk[122]) & (g21) & (!g25) & (g12) & (!g103)));
	assign g105 = (((!g24) & (!sk[123]) & (g38)) + ((g24) & (sk[123]) & (!g38)));
	assign g106 = (((!g21) & (g25) & (!sk[124]) & (!g48) & (!g105)) + ((!g21) & (!g25) & (!sk[124]) & (g48) & (!g105)) + ((!g21) & (!g25) & (!sk[124]) & (g48) & (!g105)) + ((!g21) & (!g25) & (!sk[124]) & (g48) & (!g105)));
	assign g107 = (((g35) & (!g98) & (!g102) & (!g104) & (!sk[125]) & (!g106)) + ((!g35) & (!g98) & (g102) & (!g104) & (!sk[125]) & (!g106)) + ((!g35) & (g98) & (!g102) & (g104) & (!sk[125]) & (!g106)) + ((!g35) & (!g98) & (!g102) & (g104) & (sk[125]) & (!g106)) + ((!g35) & (!g98) & (!g102) & (g104) & (sk[125]) & (!g106)));
	assign g108 = (((!g96) & (g97) & (!sk[126]) & (!g101) & (!g107)) + ((!g96) & (!g97) & (!sk[126]) & (g101) & (!g107)) + ((!g96) & (!g97) & (sk[126]) & (!g101) & (g107)));
	assign g109 = (((!sk[127]) & (g83) & (!g87) & (!g90) & (!g93) & (!g108)) + ((!sk[127]) & (!g83) & (!g87) & (g90) & (!g93) & (!g108)) + ((!sk[127]) & (!g83) & (g87) & (!g90) & (g93) & (!g108)) + ((!sk[127]) & (!g83) & (!g87) & (g90) & (g93) & (g108)));
	assign g110 = (((!i_0_) & (!i_1_) & (!sk[0]) & (i_2_)) + ((!i_0_) & (!i_1_) & (!sk[0]) & (i_2_)));
	assign g111 = (((!i_6_) & (!sk[1]) & (i_7_)) + ((!i_6_) & (!sk[1]) & (i_7_)));
	assign g112 = (((!g36) & (!g110) & (!sk[2]) & (g111)) + ((!g36) & (g110) & (!sk[2]) & (g111)));
	assign g113 = (((!i_7_) & (i_8_) & (!sk[3]) & (!g21) & (!g36)) + ((!i_7_) & (!i_8_) & (!sk[3]) & (g21) & (!g36)) + ((i_7_) & (!i_8_) & (sk[3]) & (!g21) & (!g36)) + ((!i_7_) & (!i_8_) & (sk[3]) & (!g21) & (!g36)));
	assign g114 = (((g5) & (!g36) & (!g110) & (!sk[4]) & (!g111) & (!g113)) + ((!g5) & (!g36) & (g110) & (!sk[4]) & (!g111) & (!g113)) + ((!g5) & (g36) & (!g110) & (!sk[4]) & (g111) & (!g113)) + ((!g5) & (!g36) & (!g110) & (sk[4]) & (!g111) & (!g113)) + ((!g5) & (!g36) & (!g110) & (sk[4]) & (!g111) & (!g113)) + ((!g5) & (g36) & (!g110) & (!sk[4]) & (g111) & (!g113)));
	assign g115 = (((!g47) & (!g13) & (!g15) & (!g26) & (!g112) & (g114)) + ((!g47) & (g13) & (!g15) & (!g26) & (!g112) & (!g114)) + ((!g47) & (g13) & (!g15) & (!g26) & (!g112) & (!g114)) + ((!g47) & (!g13) & (!g15) & (!g26) & (!g112) & (g114)));
	assign g116 = (((i_3_) & (!sk[6]) & (i_5_)) + ((!i_3_) & (!sk[6]) & (i_5_)));
	assign g117 = (((!sk[7]) & (!g13) & (g116)) + ((!sk[7]) & (!g13) & (g116)));
	assign g118 = (((g21) & (!g42) & (!g12) & (!sk[8]) & (!g2) & (!g59)) + ((!g21) & (!g42) & (g12) & (!sk[8]) & (!g2) & (!g59)) + ((!g21) & (g42) & (g12) & (!sk[8]) & (!g2) & (!g59)) + ((!g21) & (g42) & (!g12) & (!sk[8]) & (g2) & (!g59)) + ((!g21) & (g42) & (!g12) & (!sk[8]) & (g2) & (!g59)));
	assign g119 = (((g28) & (!g48) & (!sk[9]) & (!g26) & (!g117) & (!g118)) + ((!g28) & (!g48) & (!sk[9]) & (g26) & (!g117) & (!g118)) + ((!g28) & (g48) & (!sk[9]) & (!g26) & (g117) & (!g118)) + ((!g28) & (!g48) & (sk[9]) & (!g26) & (!g117) & (!g118)) + ((!g28) & (!g48) & (sk[9]) & (!g26) & (!g117) & (!g118)) + ((!g28) & (!g48) & (sk[9]) & (!g26) & (!g117) & (!g118)) + ((!g28) & (!g48) & (sk[9]) & (!g26) & (!g117) & (!g118)));
	assign g120 = (((!sk[10]) & (!i_3_) & (i_4_)) + ((!sk[10]) & (i_3_) & (i_4_)));
	assign g121 = (((!g28) & (!sk[11]) & (g13)) + ((g28) & (sk[11]) & (!g13)));
	assign g122 = (((g42) & (!g45) & (g6) & (!g24) & (g3) & (!g111)) + ((!g42) & (!g45) & (!g6) & (!g24) & (!g3) & (g111)));
	assign g123 = (((g50) & (!sk[13]) & (g8)) + ((!g50) & (!sk[13]) & (g8)));
	assign g124 = (((!g21) & (!g2) & (!sk[14]) & (g110)) + ((!g21) & (g2) & (!sk[14]) & (g110)));
	assign g125 = (((g12) & (!g123) & (!sk[15]) & (!g105) & (!g86) & (!g124)) + ((!g12) & (!g123) & (!sk[15]) & (g105) & (!g86) & (!g124)) + ((!g12) & (g123) & (!sk[15]) & (!g105) & (g86) & (!g124)) + ((!g12) & (!g123) & (!sk[15]) & (g105) & (!g86) & (!g124)) + ((!g12) & (!g123) & (!sk[15]) & (g105) & (!g86) & (!g124)) + ((!g12) & (!g123) & (sk[15]) & (!g105) & (!g86) & (!g124)) + ((!g12) & (!g123) & (sk[15]) & (!g105) & (!g86) & (!g124)));
	assign g126 = (((!sk[16]) & (i_3_) & (!i_4_) & (!i_5_) & (!i_0_) & (!i_1_)) + ((!sk[16]) & (!i_3_) & (!i_4_) & (i_5_) & (!i_0_) & (!i_1_)) + ((!sk[16]) & (!i_3_) & (i_4_) & (!i_5_) & (i_0_) & (!i_1_)) + ((!sk[16]) & (i_3_) & (!i_4_) & (!i_5_) & (!i_0_) & (!i_1_)) + ((!sk[16]) & (!i_3_) & (!i_4_) & (i_5_) & (!i_0_) & (i_1_)) + ((sk[16]) & (!i_3_) & (!i_4_) & (!i_5_) & (!i_0_) & (i_1_)) + ((sk[16]) & (!i_3_) & (!i_4_) & (!i_5_) & (!i_0_) & (!i_1_)));
	assign g127 = (((i_0_) & (!sk[17]) & (i_1_)) + ((!i_0_) & (!sk[17]) & (i_1_)));
	assign g128 = (((!sk[18]) & (!i_3_) & (!i_4_) & (g127)) + ((!sk[18]) & (i_3_) & (!i_4_) & (g127)));
	assign g129 = (((g42) & (!sk[19]) & (g32)) + ((!g42) & (!sk[19]) & (g32)));
	assign g130 = (((g28) & (!sk[20]) & (!g75) & (!g37) & (!g99) & (!g129)) + ((!g28) & (!sk[20]) & (!g75) & (g37) & (!g99) & (!g129)) + ((!g28) & (sk[20]) & (!g75) & (!g37) & (!g99) & (!g129)) + ((!g28) & (!sk[20]) & (!g75) & (g37) & (!g99) & (!g129)) + ((!g28) & (!sk[20]) & (g75) & (!g37) & (g99) & (!g129)) + ((!g28) & (sk[20]) & (!g75) & (!g37) & (!g99) & (!g129)));
	assign g131 = (((g120) & (!g1) & (!sk[21]) & (!g48) & (!g2) & (!g38)) + ((!g120) & (!g1) & (!sk[21]) & (g48) & (!g2) & (!g38)) + ((g120) & (!g1) & (!sk[21]) & (g48) & (!g2) & (!g38)) + ((!g120) & (g1) & (!sk[21]) & (!g48) & (g2) & (!g38)) + ((!g120) & (!g1) & (sk[21]) & (!g48) & (g2) & (!g38)));
	assign g132 = (((!sk[22]) & (g12) & (!g683) & (!g128) & (!g130) & (!g131)) + ((!sk[22]) & (!g12) & (!g683) & (g128) & (!g130) & (!g131)) + ((!sk[22]) & (!g12) & (g683) & (!g128) & (g130) & (!g131)) + ((!sk[22]) & (!g12) & (g683) & (!g128) & (g130) & (!g131)) + ((!sk[22]) & (!g12) & (g683) & (!g128) & (g130) & (!g131)));
	assign g133 = (((!sk[23]) & (!g694) & (g122) & (!g125) & (!g132)) + ((!sk[23]) & (!g694) & (!g122) & (g125) & (!g132)) + ((!sk[23]) & (g694) & (!g122) & (g125) & (g132)));
	assign g134 = (((!sk[24]) & (!i_4_) & (!i_5_) & (i_6_)) + ((sk[24]) & (!i_4_) & (!i_5_) & (!i_6_)));
	assign g135 = (((!i_3_) & (i_2_) & (!sk[25]) & (!g47) & (!g134)) + ((!i_3_) & (!i_2_) & (!sk[25]) & (g47) & (!g134)) + ((i_3_) & (i_2_) & (!sk[25]) & (g47) & (g134)));
	assign g136 = (((!i_3_) & (!i_5_) & (!i_2_) & (g35) & (!g14) & (!g64)) + ((i_3_) & (!i_5_) & (i_2_) & (!g35) & (g14) & (g64)));
	assign g137 = (((!sk[27]) & (!i_7_) & (i_8_)) + ((sk[27]) & (i_7_) & (!i_8_)));
	assign g138 = (((i_3_) & (!sk[28]) & (!i_0_) & (!i_1_) & (!g137) & (!g85)) + ((!i_3_) & (!sk[28]) & (!i_0_) & (i_1_) & (!g137) & (!g85)) + ((!i_3_) & (!sk[28]) & (i_0_) & (!i_1_) & (g137) & (!g85)) + ((!i_3_) & (!sk[28]) & (!i_0_) & (i_1_) & (g137) & (g85)));
	assign g139 = (((!i_3_) & (i_5_) & (!g28) & (!sk[29]) & (!g24)) + ((!i_3_) & (!i_5_) & (g28) & (!sk[29]) & (!g24)) + ((!i_3_) & (i_5_) & (g28) & (!sk[29]) & (!g24)));
	assign g140 = (((g27) & (!g6) & (!sk[30]) & (!g36) & (!g138) & (!g139)) + ((!g27) & (!g6) & (!sk[30]) & (g36) & (!g138) & (!g139)) + ((!g27) & (g6) & (!sk[30]) & (!g36) & (g138) & (!g139)) + ((g27) & (!g6) & (!sk[30]) & (!g36) & (!g138) & (!g139)) + ((!g27) & (!g6) & (!sk[30]) & (g36) & (!g138) & (!g139)) + ((!g27) & (!g6) & (sk[30]) & (!g36) & (!g138) & (!g139)));
	assign g141 = (((!g35) & (!sk[31]) & (g24)) + ((g35) & (sk[31]) & (!g24)));
	assign g142 = (((i_3_) & (!g42) & (!g8) & (!sk[32]) & (!g45) & (!g141)) + ((!i_3_) & (!g42) & (g8) & (!sk[32]) & (!g45) & (!g141)) + ((!i_3_) & (g42) & (g8) & (!sk[32]) & (!g45) & (!g141)) + ((!i_3_) & (g42) & (!g8) & (!sk[32]) & (g45) & (!g141)) + ((!i_3_) & (!g42) & (!g8) & (sk[32]) & (!g45) & (g141)));
	assign g143 = (((!i_8_) & (g51) & (!g64) & (!sk[33]) & (!g142)) + ((!i_8_) & (!g51) & (g64) & (!sk[33]) & (!g142)) + ((i_8_) & (!g51) & (!g64) & (sk[33]) & (!g142)) + ((!i_8_) & (!g51) & (!g64) & (sk[33]) & (!g142)) + ((!i_8_) & (!g51) & (!g64) & (sk[33]) & (!g142)));
	assign g144 = (((!sk[34]) & (i_1_) & (!g135) & (!g136) & (!g140) & (!g143)) + ((!sk[34]) & (!i_1_) & (!g135) & (g136) & (!g140) & (!g143)) + ((!sk[34]) & (!i_1_) & (g135) & (!g136) & (g140) & (!g143)) + ((sk[34]) & (!i_1_) & (!g135) & (!g136) & (g140) & (g143)) + ((sk[34]) & (!i_1_) & (!g135) & (!g136) & (g140) & (g143)));
	assign g145 = (((i_6_) & (!sk[35]) & (!g137) & (!g51) & (!g33) & (!g85)) + ((!i_6_) & (!sk[35]) & (!g137) & (g51) & (!g33) & (!g85)) + ((!i_6_) & (!sk[35]) & (g137) & (!g51) & (g33) & (!g85)) + ((!i_6_) & (!sk[35]) & (g137) & (g51) & (!g33) & (g85)));
	assign g146 = (((g27) & (!sk[36]) & (!i_6_) & (!g47) & (!g24) & (!g3)) + ((!g27) & (!sk[36]) & (!i_6_) & (g47) & (!g24) & (!g3)) + ((!g27) & (!sk[36]) & (i_6_) & (!g47) & (g24) & (!g3)) + ((!g27) & (!sk[36]) & (!i_6_) & (g47) & (!g24) & (g3)) + ((!g27) & (!sk[36]) & (i_6_) & (g47) & (!g24) & (g3)));
	assign g147 = (((g37) & (!sk[37]) & (!g38) & (!g110) & (!g145) & (!g146)) + ((!g37) & (!sk[37]) & (!g38) & (g110) & (!g145) & (!g146)) + ((!g37) & (!sk[37]) & (g38) & (!g110) & (g145) & (!g146)) + ((!g37) & (sk[37]) & (!g38) & (!g110) & (!g145) & (!g146)) + ((!g37) & (sk[37]) & (g38) & (!g110) & (!g145) & (!g146)) + ((!g37) & (sk[37]) & (!g38) & (!g110) & (!g145) & (!g146)));
	assign g148 = (((g11) & (!g42) & (!sk[38]) & (!g47) & (!g64) & (!g111)) + ((!g11) & (!g42) & (!sk[38]) & (g47) & (!g64) & (!g111)) + ((!g11) & (g42) & (!sk[38]) & (!g47) & (g64) & (!g111)) + ((!g11) & (g42) & (!sk[38]) & (g47) & (g64) & (!g111)) + ((!g11) & (g42) & (sk[38]) & (!g47) & (!g64) & (g111)));
	assign g149 = (((!g21) & (!sk[39]) & (g23) & (!g7) & (!g100)) + ((!g21) & (!sk[39]) & (!g23) & (g7) & (!g100)) + ((!g21) & (!sk[39]) & (!g23) & (g7) & (!g100)) + ((!g21) & (sk[39]) & (!g23) & (!g7) & (g100)));
	assign g150 = (((!sk[40]) & (!g12) & (!g59) & (g13)) + ((sk[40]) & (g12) & (!g59) & (!g13)));
	assign g151 = (((!g25) & (g12) & (!sk[41]) & (!g3) & (!g150)) + ((!g25) & (!g12) & (!sk[41]) & (g3) & (!g150)) + ((g25) & (!g12) & (sk[41]) & (!g3) & (!g150)) + ((!g25) & (!g12) & (sk[41]) & (!g3) & (!g150)) + ((!g25) & (!g12) & (sk[41]) & (!g3) & (!g150)));
	assign g152 = (((!sk[42]) & (g6) & (!g77) & (!g148) & (!g149) & (!g151)) + ((!sk[42]) & (!g6) & (!g77) & (g148) & (!g149) & (!g151)) + ((!sk[42]) & (!g6) & (g77) & (!g148) & (g149) & (!g151)) + ((sk[42]) & (!g6) & (!g77) & (!g148) & (!g149) & (g151)) + ((!sk[42]) & (g6) & (!g77) & (!g148) & (!g149) & (g151)));
	assign g153 = (((!sk[43]) & (!g670) & (!g147) & (g152)) + ((!sk[43]) & (g670) & (g147) & (g152)));
	assign g154 = (((g115) & (!g119) & (!g133) & (!g144) & (!sk[44]) & (!g153)) + ((!g115) & (!g119) & (g133) & (!g144) & (!sk[44]) & (!g153)) + ((!g115) & (g119) & (!g133) & (g144) & (!sk[44]) & (!g153)) + ((g115) & (g119) & (g133) & (g144) & (!sk[44]) & (g153)));
	assign g155 = (((!g11) & (!g27) & (!sk[45]) & (g28)) + ((!g11) & (!g27) & (!sk[45]) & (g28)));
	assign g156 = (((!g23) & (!g36) & (g7) & (!sk[46]) & (!g129)) + ((!g23) & (g36) & (!g7) & (!sk[46]) & (!g129)) + ((!g23) & (!g36) & (!g7) & (sk[46]) & (g129)));
	assign g157 = (((!sk[47]) & (!g47) & (g75) & (!g155) & (!g156)) + ((!sk[47]) & (!g47) & (!g75) & (g155) & (!g156)) + ((sk[47]) & (!g47) & (!g75) & (!g155) & (!g156)) + ((!sk[47]) & (!g47) & (g75) & (!g155) & (!g156)));
	assign g158 = (((!g1) & (!sk[48]) & (g59)) + ((!g1) & (sk[48]) & (!g59)));
	assign g159 = (((!sk[49]) & (!g21) & (g48)) + ((!sk[49]) & (!g21) & (g48)));
	assign g160 = (((!sk[50]) & (!g42) & (g12) & (!g84) & (!g159)) + ((!sk[50]) & (!g42) & (!g12) & (g84) & (!g159)) + ((!sk[50]) & (!g42) & (g12) & (g84) & (!g159)) + ((sk[50]) & (g42) & (!g12) & (!g84) & (g159)));
	assign g161 = (((!sk[51]) & (!g11) & (g110)) + ((!sk[51]) & (!g11) & (g110)));
	assign g162 = (((g28) & (!g2) & (!sk[52]) & (!g24) & (!g32) & (!g161)) + ((!g28) & (!g2) & (!sk[52]) & (g24) & (!g32) & (!g161)) + ((g28) & (!g2) & (!sk[52]) & (!g24) & (!g32) & (g161)) + ((!g28) & (g2) & (!sk[52]) & (!g24) & (g32) & (!g161)));
	assign g163 = (((i_7_) & (!i_8_) & (!g45) & (!sk[53]) & (!g13) & (!g88)) + ((!i_7_) & (!i_8_) & (g45) & (!sk[53]) & (!g13) & (!g88)) + ((!i_7_) & (i_8_) & (!g45) & (!sk[53]) & (g13) & (!g88)) + ((i_7_) & (i_8_) & (!g45) & (!sk[53]) & (!g13) & (g88)) + ((i_7_) & (!i_8_) & (!g45) & (!sk[53]) & (!g13) & (!g88)));
	assign g164 = (((!sk[54]) & (g2) & (!g158) & (!g160) & (!g162) & (!g163)) + ((!sk[54]) & (!g2) & (!g158) & (g160) & (!g162) & (!g163)) + ((!sk[54]) & (!g2) & (g158) & (!g160) & (g162) & (!g163)) + ((sk[54]) & (!g2) & (!g158) & (!g160) & (!g162) & (!g163)) + ((!sk[54]) & (g2) & (!g158) & (!g160) & (!g162) & (!g163)));
	assign g165 = (((!g27) & (!sk[55]) & (!g59) & (g60)) + ((!g27) & (!sk[55]) & (!g59) & (g60)));
	assign g166 = (((!sk[56]) & (!i_5_) & (g42) & (!g2) & (!g165)) + ((!sk[56]) & (!i_5_) & (!g42) & (g2) & (!g165)) + ((sk[56]) & (i_5_) & (!g42) & (!g2) & (!g165)) + ((sk[56]) & (!i_5_) & (!g42) & (!g2) & (!g165)) + ((sk[56]) & (!i_5_) & (!g42) & (!g2) & (!g165)));
	assign g167 = (((!sk[57]) & (!g14) & (g134)) + ((!sk[57]) & (g14) & (g134)));
	assign g168 = (((!i_0_) & (!i_2_) & (g35) & (g75) & (!sk[58]) & (!g167)) + ((i_0_) & (!i_2_) & (!g35) & (!g75) & (!sk[58]) & (!g167)) + ((!i_0_) & (!i_2_) & (g35) & (!g75) & (!sk[58]) & (!g167)) + ((!i_0_) & (i_2_) & (!g35) & (g75) & (!sk[58]) & (!g167)) + ((i_0_) & (i_2_) & (!g35) & (!g75) & (!sk[58]) & (g167)));
	assign g169 = (((!g50) & (!sk[59]) & (i_6_) & (!g42) & (!g47)) + ((!g50) & (!sk[59]) & (!i_6_) & (g42) & (!g47)) + ((g50) & (!sk[59]) & (i_6_) & (g42) & (g47)));
	assign g170 = (((!sk[60]) & (!i_3_) & (i_5_) & (!g25) & (!g12)) + ((!sk[60]) & (!i_3_) & (!i_5_) & (g25) & (!g12)) + ((sk[60]) & (i_3_) & (!i_5_) & (!g25) & (g12)));
	assign g171 = (((!i_3_) & (!sk[61]) & (i_5_) & (!g2) & (!g13)) + ((!i_3_) & (!sk[61]) & (!i_5_) & (g2) & (!g13)) + ((!i_3_) & (!sk[61]) & (i_5_) & (g2) & (!g13)));
	assign g172 = (((!g32) & (!sk[62]) & (g121) & (!g170) & (!g171)) + ((!g32) & (!sk[62]) & (!g121) & (g170) & (!g171)) + ((!g32) & (sk[62]) & (!g121) & (!g170) & (!g171)) + ((!g32) & (!sk[62]) & (g121) & (!g170) & (!g171)));
	assign g173 = (((g127) & (!i_2_) & (!sk[63]) & (!g8) & (!g45) & (!g12)) + ((!g127) & (!i_2_) & (!sk[63]) & (g8) & (!g45) & (!g12)) + ((!g127) & (i_2_) & (!sk[63]) & (!g8) & (g45) & (!g12)) + ((g127) & (!i_2_) & (!sk[63]) & (g8) & (!g45) & (!g12)) + ((g127) & (i_2_) & (!sk[63]) & (!g8) & (!g45) & (g12)));
	assign g174 = (((!g11) & (g8) & (!sk[64]) & (!g29) & (!g91)) + ((!g11) & (!g8) & (!sk[64]) & (g29) & (!g91)) + ((!g11) & (!g8) & (!sk[64]) & (g29) & (!g91)) + ((!g11) & (g8) & (!sk[64]) & (!g29) & (g91)));
	assign g175 = (((!sk[65]) & (!g25) & (g45) & (!g22) & (!g6)) + ((!sk[65]) & (!g25) & (!g45) & (g22) & (!g6)) + ((!sk[65]) & (!g25) & (!g45) & (g22) & (!g6)) + ((sk[65]) & (!g25) & (!g45) & (!g22) & (g6)));
	assign g176 = (((g28) & (!g25) & (!g59) & (!g7) & (!sk[66]) & (!g110)) + ((!g28) & (!g25) & (g59) & (!g7) & (!sk[66]) & (!g110)) + ((g28) & (!g25) & (!g59) & (!g7) & (!sk[66]) & (!g110)) + ((!g28) & (!g25) & (!g59) & (g7) & (sk[66]) & (!g110)) + ((g28) & (!g25) & (!g59) & (!g7) & (!sk[66]) & (g110)) + ((!g28) & (g25) & (!g59) & (g7) & (!sk[66]) & (!g110)));
	assign g177 = (((!g173) & (!sk[67]) & (g174) & (!g175) & (!g176)) + ((!g173) & (!sk[67]) & (!g174) & (g175) & (!g176)) + ((!g173) & (sk[67]) & (!g174) & (!g175) & (!g176)));
	assign g178 = (((g11) & (!g9) & (!sk[68]) & (!g169) & (!g172) & (!g177)) + ((!g11) & (!g9) & (!sk[68]) & (g169) & (!g172) & (!g177)) + ((!g11) & (g9) & (!sk[68]) & (!g169) & (g172) & (!g177)) + ((g11) & (!g9) & (!sk[68]) & (!g169) & (g172) & (g177)) + ((!g11) & (!g9) & (sk[68]) & (!g169) & (g172) & (g177)));
	assign g179 = (((g35) & (!sk[69]) & (!g21) & (!g12) & (!g24) & (!g26)) + ((!g35) & (!sk[69]) & (!g21) & (g12) & (!g24) & (!g26)) + ((g35) & (!sk[69]) & (!g21) & (!g12) & (!g24) & (g26)) + ((!g35) & (!sk[69]) & (g21) & (!g12) & (g24) & (!g26)) + ((!g35) & (!sk[69]) & (!g21) & (g12) & (!g24) & (!g26)));
	assign g180 = (((!i_3_) & (!i_4_) & (i_5_) & (!g127) & (g63) & (g51)) + ((i_3_) & (i_4_) & (i_5_) & (g127) & (g63) & (!g51)));
	assign g181 = (((!sk[71]) & (!g45) & (g110)) + ((!sk[71]) & (!g45) & (g110)));
	assign g182 = (((!i_6_) & (i_7_) & (!i_8_) & (g75) & (!g181) & (!g105)) + ((i_6_) & (i_7_) & (i_8_) & (!g75) & (g181) & (!g105)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g75) & (!g181) & (!g105)));
	assign g183 = (((!sk[73]) & (i_3_) & (!i_5_) & (!g127) & (!g28) & (!g123)) + ((!sk[73]) & (!i_3_) & (!i_5_) & (g127) & (!g28) & (!g123)) + ((!sk[73]) & (!i_3_) & (i_5_) & (!g127) & (g28) & (!g123)) + ((!sk[73]) & (!i_3_) & (!i_5_) & (g127) & (!g28) & (g123)) + ((!sk[73]) & (i_3_) & (i_5_) & (g127) & (g28) & (!g123)));
	assign g184 = (((!g59) & (!sk[74]) & (g110)) + ((!g59) & (!sk[74]) & (g110)));
	assign g185 = (((!sk[75]) & (!g2) & (g23) & (!g70) & (!g184)) + ((!sk[75]) & (!g2) & (!g23) & (g70) & (!g184)) + ((!sk[75]) & (g2) & (!g23) & (g70) & (!g184)) + ((sk[75]) & (!g2) & (!g23) & (!g70) & (g184)));
	assign g186 = (((!sk[76]) & (g45) & (!g48) & (!g2) & (!g24) & (!g184)) + ((!sk[76]) & (!g45) & (!g48) & (g2) & (!g24) & (!g184)) + ((!sk[76]) & (!g45) & (!g48) & (g2) & (!g24) & (g184)) + ((!sk[76]) & (!g45) & (g48) & (!g2) & (g24) & (!g184)) + ((sk[76]) & (!g45) & (g48) & (!g2) & (!g24) & (!g184)));
	assign g187 = (((!i_3_) & (!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (!i_8_)));
	assign g188 = (((!sk[78]) & (!i_3_) & (i_5_) & (!g35) & (!g42)) + ((!sk[78]) & (!i_3_) & (!i_5_) & (g35) & (!g42)) + ((!sk[78]) & (i_3_) & (!i_5_) & (g35) & (g42)));
	assign g189 = (((!sk[79]) & (!g3) & (g110)) + ((!sk[79]) & (g3) & (g110)));
	assign g190 = (((!i_6_) & (!sk[80]) & (!g63) & (g188) & (!g181) & (!g189)) + ((!i_6_) & (sk[80]) & (!g63) & (!g188) & (!g181) & (!g189)) + ((!i_6_) & (!sk[80]) & (g63) & (!g188) & (g181) & (!g189)) + ((i_6_) & (!sk[80]) & (!g63) & (!g188) & (!g181) & (!g189)) + ((i_6_) & (!sk[80]) & (!g63) & (!g188) & (!g181) & (!g189)) + ((!i_6_) & (sk[80]) & (!g63) & (!g188) & (!g181) & (!g189)));
	assign g191 = (((!sk[81]) & (!g185) & (g186) & (!g657) & (!g190)) + ((!sk[81]) & (!g185) & (!g186) & (g657) & (!g190)) + ((!sk[81]) & (!g185) & (!g186) & (g657) & (g190)));
	assign g192 = (((!sk[82]) & (g179) & (!g180) & (!g182) & (!g183) & (!g191)) + ((!sk[82]) & (!g179) & (!g180) & (g182) & (!g183) & (!g191)) + ((!sk[82]) & (!g179) & (g180) & (!g182) & (g183) & (!g191)) + ((sk[82]) & (!g179) & (!g180) & (!g182) & (!g183) & (g191)));
	assign g193 = (((!g23) & (g3) & (!sk[83]) & (!g7) & (!g181)) + ((!g23) & (g3) & (!sk[83]) & (g7) & (!g181)) + ((!g23) & (!g3) & (!sk[83]) & (g7) & (!g181)) + ((!g23) & (!g3) & (sk[83]) & (!g7) & (g181)));
	assign g194 = (((!sk[84]) & (!g21) & (g6)) + ((!sk[84]) & (!g21) & (g6)));
	assign g195 = (((!g8) & (g13) & (!sk[85]) & (!g181) & (!g194)) + ((g8) & (!g13) & (!sk[85]) & (g181) & (!g194)) + ((!g8) & (!g13) & (!sk[85]) & (g181) & (!g194)) + ((!g8) & (!g13) & (sk[85]) & (!g181) & (g194)));
	assign g196 = (((g27) & (!g23) & (!g3) & (!g110) & (!sk[86]) & (!g194)) + ((!g27) & (!g23) & (g3) & (!g110) & (!sk[86]) & (!g194)) + ((!g27) & (!g23) & (g3) & (!g110) & (!sk[86]) & (!g194)) + ((!g27) & (g23) & (!g3) & (g110) & (!sk[86]) & (!g194)) + ((!g27) & (!g23) & (!g3) & (g110) & (sk[86]) & (g194)));
	assign g197 = (((g47) & (!g73) & (!g193) & (!g195) & (!sk[87]) & (!g196)) + ((!g47) & (!g73) & (g193) & (!g195) & (!sk[87]) & (!g196)) + ((!g47) & (g73) & (!g193) & (g195) & (!sk[87]) & (!g196)) + ((!g47) & (!g73) & (!g193) & (!g195) & (sk[87]) & (!g196)) + ((!g47) & (!g73) & (!g193) & (!g195) & (sk[87]) & (!g196)));
	assign g198 = (((!sk[88]) & (g166) & (!g168) & (!g178) & (!g192) & (!g197)) + ((!sk[88]) & (!g166) & (!g168) & (g178) & (!g192) & (!g197)) + ((!sk[88]) & (!g166) & (g168) & (!g178) & (g192) & (!g197)) + ((!sk[88]) & (g166) & (!g168) & (g178) & (g192) & (g197)));
	assign g199 = (((!sk[89]) & (g109) & (!g154) & (!g157) & (!g164) & (!g198)) + ((!sk[89]) & (!g109) & (!g154) & (g157) & (!g164) & (!g198)) + ((!sk[89]) & (!g109) & (g154) & (!g157) & (g164) & (!g198)) + ((!sk[89]) & (g109) & (g154) & (g157) & (g164) & (g198)));
	assign g200 = (((!sk[90]) & (g27) & (!g45) & (!g23) & (!g36) & (!g121)) + ((!sk[90]) & (!g27) & (!g45) & (g23) & (!g36) & (!g121)) + ((!sk[90]) & (!g27) & (g45) & (!g23) & (g36) & (!g121)) + ((sk[90]) & (!g27) & (!g45) & (!g23) & (!g36) & (g121)) + ((sk[90]) & (!g27) & (!g45) & (!g23) & (!g36) & (!g121)));
	assign g201 = (((g50) & (!i_6_) & (!g137) & (!g94) & (!sk[91]) & (!g88)) + ((!g50) & (!i_6_) & (g137) & (!g94) & (!sk[91]) & (!g88)) + ((!g50) & (i_6_) & (!g137) & (g94) & (!sk[91]) & (!g88)) + ((!g50) & (!i_6_) & (g137) & (!g94) & (!sk[91]) & (g88)) + ((g50) & (i_6_) & (g137) & (g94) & (!sk[91]) & (!g88)));
	assign g202 = (((!g45) & (!sk[92]) & (g37) & (!g13) & (!g201)) + ((!g45) & (!sk[92]) & (!g37) & (g13) & (!g201)) + ((!g45) & (!sk[92]) & (!g37) & (g13) & (!g201)) + ((!g45) & (sk[92]) & (!g37) & (!g13) & (!g201)) + ((g45) & (!sk[92]) & (g37) & (!g13) & (!g201)));
	assign g203 = (((!sk[93]) & (i_6_) & (!g63) & (!g21) & (!g13) & (!g84)) + ((!sk[93]) & (!i_6_) & (!g63) & (g21) & (!g13) & (!g84)) + ((!sk[93]) & (!i_6_) & (g63) & (!g21) & (g13) & (!g84)) + ((!sk[93]) & (i_6_) & (g63) & (!g21) & (!g13) & (g84)) + ((sk[93]) & (!i_6_) & (g63) & (!g21) & (!g13) & (!g84)));
	assign g204 = (((!sk[94]) & (i_6_) & (!i_8_) & (!g32) & (!g105) & (!g141)) + ((!sk[94]) & (!i_6_) & (!i_8_) & (g32) & (!g105) & (!g141)) + ((!sk[94]) & (!i_6_) & (!i_8_) & (g32) & (!g105) & (g141)) + ((!sk[94]) & (!i_6_) & (i_8_) & (!g32) & (g105) & (!g141)) + ((!sk[94]) & (i_6_) & (i_8_) & (!g32) & (!g105) & (!g141)));
	assign g205 = (((!g23) & (!sk[95]) & (!g70) & (g204)) + ((g23) & (sk[95]) & (!g70) & (!g204)) + ((!g23) & (sk[95]) & (!g70) & (!g204)));
	assign g206 = (((!sk[96]) & (g150) & (!g200) & (!g202) & (!g203) & (!g205)) + ((!sk[96]) & (!g150) & (!g200) & (g202) & (!g203) & (!g205)) + ((!sk[96]) & (!g150) & (g200) & (!g202) & (g203) & (!g205)) + ((!sk[96]) & (!g150) & (!g200) & (g202) & (!g203) & (g205)));
	assign g207 = (((!i_3_) & (!sk[97]) & (i_5_) & (!g8) & (!g24)) + ((!i_3_) & (!sk[97]) & (!i_5_) & (g8) & (!g24)) + ((!i_3_) & (!sk[97]) & (!i_5_) & (g8) & (!g24)));
	assign g208 = (((i_6_) & (!g42) & (!g46) & (!sk[98]) & (!g47) & (!g38)) + ((!i_6_) & (!g42) & (g46) & (!sk[98]) & (!g47) & (!g38)) + ((!i_6_) & (!g42) & (g46) & (!sk[98]) & (g47) & (!g38)) + ((!i_6_) & (g42) & (!g46) & (!sk[98]) & (g47) & (!g38)) + ((i_6_) & (g42) & (!g46) & (!sk[98]) & (g47) & (!g38)));
	assign g209 = (((g127) & (!sk[99]) & (!i_2_) & (!g8) & (!g22) & (!g59)) + ((!g127) & (!sk[99]) & (!i_2_) & (g8) & (!g22) & (!g59)) + ((!g127) & (!sk[99]) & (i_2_) & (!g8) & (g22) & (!g59)) + ((g127) & (!sk[99]) & (!i_2_) & (!g8) & (g22) & (!g59)) + ((g127) & (!sk[99]) & (i_2_) & (g8) & (!g22) & (!g59)));
	assign g210 = (((g28) & (!g26) & (!sk[100]) & (!g208) & (!g644) & (!g209)) + ((!g28) & (!g26) & (!sk[100]) & (g208) & (!g644) & (!g209)) + ((!g28) & (g26) & (!sk[100]) & (!g208) & (g644) & (!g209)) + ((!g28) & (!g26) & (sk[100]) & (!g208) & (g644) & (!g209)) + ((!g28) & (!g26) & (sk[100]) & (!g208) & (g644) & (!g209)));
	assign g211 = (((g1) & (!g47) & (!g64) & (!sk[101]) & (!g207) & (!g210)) + ((!g1) & (!g47) & (g64) & (!sk[101]) & (!g207) & (!g210)) + ((!g1) & (g47) & (!g64) & (!sk[101]) & (g207) & (!g210)) + ((g1) & (!g47) & (!g64) & (!sk[101]) & (!g207) & (g210)) + ((!g1) & (!g47) & (!g64) & (sk[101]) & (!g207) & (g210)) + ((!g1) & (!g47) & (!g64) & (sk[101]) & (!g207) & (g210)));
	assign g212 = (((!g45) & (!g23) & (!sk[102]) & (g24)) + ((!g45) & (!g23) & (sk[102]) & (!g24)));
	assign g213 = (((!sk[103]) & (!g50) & (i_6_) & (!g42) & (!g137)) + ((!sk[103]) & (!g50) & (!i_6_) & (g42) & (!g137)) + ((!sk[103]) & (g50) & (i_6_) & (g42) & (g137)));
	assign g214 = (((g2) & (!g73) & (!sk[104]) & (!g38) & (!g29) & (!g213)) + ((!g2) & (!g73) & (!sk[104]) & (g38) & (!g29) & (!g213)) + ((!g2) & (g73) & (!sk[104]) & (!g38) & (g29) & (!g213)) + ((!g2) & (!g73) & (!sk[104]) & (g38) & (!g29) & (!g213)) + ((!g2) & (!g73) & (!sk[104]) & (g38) & (!g29) & (!g213)) + ((!g2) & (!g73) & (sk[104]) & (!g38) & (!g29) & (!g213)) + ((!g2) & (!g73) & (sk[104]) & (!g38) & (!g29) & (!g213)));
	assign g215 = (((i_4_) & (!i_5_) & (!g6) & (!sk[105]) & (!g13) & (!g214)) + ((!i_4_) & (!i_5_) & (g6) & (!sk[105]) & (!g13) & (!g214)) + ((!i_4_) & (i_5_) & (!g6) & (!sk[105]) & (g13) & (!g214)) + ((!i_4_) & (!i_5_) & (!g6) & (sk[105]) & (!g13) & (g214)) + ((!i_4_) & (!i_5_) & (!g6) & (sk[105]) & (!g13) & (g214)) + ((!i_4_) & (!i_5_) & (!g6) & (sk[105]) & (!g13) & (g214)) + ((!i_4_) & (!i_5_) & (!g6) & (sk[105]) & (g13) & (g214)));
	assign g216 = (((!i_1_) & (!sk[106]) & (g135) & (!g212) & (!g215)) + ((!i_1_) & (!sk[106]) & (!g135) & (g212) & (!g215)) + ((!i_1_) & (sk[106]) & (!g135) & (!g212) & (g215)) + ((i_1_) & (!sk[106]) & (g135) & (!g212) & (g215)));
	assign g217 = (((!sk[107]) & (!i_3_) & (!i_5_) & (i_6_)) + ((sk[107]) & (!i_3_) & (i_5_) & (!i_6_)));
	assign g218 = (((g42) & (!sk[108]) & (g217)) + ((!g42) & (!sk[108]) & (g217)));
	assign g219 = (((g63) & (!sk[109]) & (g15)) + ((!g63) & (!sk[109]) & (g15)));
	assign g220 = (((!sk[110]) & (!i_3_) & (i_1_) & (!i_2_) & (!g219)) + ((!sk[110]) & (!i_3_) & (!i_1_) & (i_2_) & (!g219)) + ((!sk[110]) & (!i_3_) & (i_1_) & (!i_2_) & (g219)));
	assign g221 = (((g27) & (!g35) & (!sk[111]) & (!g28) & (!g1) & (!g36)) + ((!g27) & (!g35) & (!sk[111]) & (g28) & (!g1) & (!g36)) + ((!g27) & (g35) & (!sk[111]) & (!g28) & (g1) & (!g36)) + ((!g27) & (!g35) & (!sk[111]) & (g28) & (!g1) & (!g36)) + ((!g27) & (g35) & (sk[111]) & (!g28) & (!g1) & (!g36)));
	assign g222 = (((!sk[112]) & (g23) & (!g59) & (!g13) & (!g105) & (!g221)) + ((!sk[112]) & (!g23) & (!g59) & (g13) & (!g105) & (!g221)) + ((!sk[112]) & (g23) & (!g59) & (!g13) & (!g105) & (!g221)) + ((!sk[112]) & (!g23) & (g59) & (!g13) & (g105) & (!g221)) + ((!sk[112]) & (!g23) & (g59) & (!g13) & (g105) & (!g221)) + ((!sk[112]) & (!g23) & (!g59) & (g13) & (g105) & (!g221)));
	assign g223 = (((!g27) & (!sk[113]) & (g43) & (!g23) & (!g3)) + ((!g27) & (!sk[113]) & (!g43) & (g23) & (!g3)) + ((g27) & (sk[113]) & (!g43) & (!g23) & (!g3)) + ((!g27) & (sk[113]) & (!g43) & (!g23) & (!g3)));
	assign g224 = (((i_7_) & (!g218) & (!g220) & (!g222) & (!sk[114]) & (!g223)) + ((!i_7_) & (!g218) & (g220) & (!g222) & (!sk[114]) & (!g223)) + ((!i_7_) & (g218) & (!g220) & (g222) & (!sk[114]) & (!g223)) + ((i_7_) & (!g218) & (!g220) & (g222) & (!sk[114]) & (g223)) + ((!i_7_) & (!g218) & (!g220) & (g222) & (sk[114]) & (g223)));
	assign g225 = (((!sk[115]) & (!i_3_) & (!i_4_) & (i_6_)) + ((sk[115]) & (!i_3_) & (!i_4_) & (!i_6_)));
	assign g226 = (((g63) & (!g41) & (!g1) & (!g36) & (!sk[116]) & (!g225)) + ((!g63) & (!g41) & (g1) & (!g36) & (!sk[116]) & (!g225)) + ((!g63) & (g41) & (!g1) & (!g36) & (sk[116]) & (!g225)) + ((!g63) & (g41) & (!g1) & (g36) & (!sk[116]) & (!g225)) + ((g63) & (!g41) & (!g1) & (!g36) & (!sk[116]) & (g225)));
	assign g227 = (((i_6_) & (!i_7_) & (!i_8_) & (!g100) & (!sk[117]) & (!g129)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g100) & (!sk[117]) & (!g129)) + ((!i_6_) & (i_7_) & (!i_8_) & (g100) & (!sk[117]) & (!g129)) + ((!i_6_) & (!i_7_) & (i_8_) & (g100) & (!sk[117]) & (!g129)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g100) & (sk[117]) & (g129)));
	assign g228 = (((!g186) & (!sk[118]) & (!g226) & (g227)) + ((!g186) & (sk[118]) & (!g226) & (!g227)));
	assign g229 = (((!g23) & (!g71) & (!sk[119]) & (g161)) + ((!g23) & (!g71) & (!sk[119]) & (g161)) + ((!g23) & (g71) & (sk[119]) & (!g161)));
	assign g230 = (((!i_3_) & (!sk[120]) & (!i_1_) & (i_2_)) + ((!i_3_) & (!sk[120]) & (i_1_) & (i_2_)));
	assign g231 = (((g50) & (!g8) & (!g12) & (!sk[121]) & (!g57) & (!g230)) + ((!g50) & (!g8) & (g12) & (!sk[121]) & (!g57) & (!g230)) + ((g50) & (g8) & (!g12) & (!sk[121]) & (g57) & (!g230)) + ((!g50) & (g8) & (!g12) & (!sk[121]) & (g57) & (!g230)) + ((g50) & (!g8) & (g12) & (!sk[121]) & (!g57) & (g230)));
	assign g232 = (((!i_6_) & (!i_7_) & (i_8_) & (!g75) & (!g158) & (!g231)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g75) & (!g158) & (!g231)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g75) & (!g158) & (!g231)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g75) & (!g158) & (!g231)) + ((i_6_) & (i_7_) & (!i_8_) & (!g75) & (!g158) & (!g231)) + ((!i_6_) & (!i_7_) & (!i_8_) & (!g75) & (!g158) & (!g231)));
	assign g233 = (((g25) & (!g194) & (!sk[123]) & (!g229) & (!g631) & (!g232)) + ((!g25) & (!g194) & (!sk[123]) & (g229) & (!g631) & (!g232)) + ((!g25) & (g194) & (!sk[123]) & (!g229) & (g631) & (!g232)) + ((g25) & (!g194) & (!sk[123]) & (!g229) & (g631) & (g232)) + ((!g25) & (!g194) & (sk[123]) & (!g229) & (g631) & (g232)));
	assign g234 = (((g30) & (!g216) & (!g224) & (!g228) & (!sk[124]) & (!g233)) + ((!g30) & (!g216) & (g224) & (!g228) & (!sk[124]) & (!g233)) + ((!g30) & (g216) & (!g224) & (g228) & (!sk[124]) & (!g233)) + ((!g30) & (g216) & (g224) & (g228) & (!sk[124]) & (g233)));
	assign g235 = (((g35) & (!g21) & (!g8) & (!sk[125]) & (!g25) & (!g32)) + ((!g35) & (!g21) & (g8) & (!sk[125]) & (!g25) & (!g32)) + ((!g35) & (g21) & (!g8) & (!sk[125]) & (g25) & (!g32)) + ((g35) & (!g21) & (!g8) & (!sk[125]) & (!g25) & (!g32)) + ((!g35) & (!g21) & (g8) & (!sk[125]) & (!g25) & (g32)));
	assign g236 = (((g6) & (!sk[126]) & (!g73) & (!g49) & (!g60) & (!g235)) + ((!g6) & (!sk[126]) & (!g73) & (g49) & (!g60) & (!g235)) + ((!g6) & (!sk[126]) & (g73) & (!g49) & (g60) & (!g235)) + ((!g6) & (sk[126]) & (!g73) & (!g49) & (!g60) & (!g235)) + ((!g6) & (sk[126]) & (!g73) & (!g49) & (!g60) & (!g235)) + ((!g6) & (sk[126]) & (!g73) & (!g49) & (!g60) & (!g235)) + ((!g6) & (!sk[126]) & (!g73) & (g49) & (!g60) & (!g235)));
	assign g237 = (((!sk[127]) & (!g21) & (g8) & (!g24) & (!g69)) + ((!sk[127]) & (!g21) & (!g8) & (g24) & (!g69)) + ((!sk[127]) & (!g21) & (!g8) & (g24) & (g69)) + ((sk[127]) & (!g21) & (!g8) & (!g24) & (g69)) + ((!sk[127]) & (g21) & (g8) & (!g24) & (g69)));
	assign g238 = (((!sk[0]) & (g11) & (!g1) & (!g23) & (!g3) & (!g141)) + ((!sk[0]) & (!g11) & (!g1) & (g23) & (!g3) & (!g141)) + ((!sk[0]) & (!g11) & (g1) & (!g23) & (g3) & (!g141)) + ((sk[0]) & (!g11) & (!g1) & (!g23) & (!g3) & (g141)) + ((sk[0]) & (!g11) & (!g1) & (!g23) & (g3) & (!g141)));
	assign g239 = (((g11) & (!sk[1]) & (!g45) & (!g2) & (!g23) & (!g13)) + ((!g11) & (!sk[1]) & (!g45) & (g2) & (!g23) & (!g13)) + ((!g11) & (!sk[1]) & (g45) & (!g2) & (g23) & (!g13)) + ((!g11) & (!sk[1]) & (!g45) & (g2) & (!g23) & (!g13)) + ((!g11) & (sk[1]) & (!g45) & (!g2) & (!g23) & (!g13)));
	assign g240 = (((!g25) & (g120) & (!g12) & (!sk[2]) & (!g181)) + ((!g25) & (!g120) & (g12) & (!sk[2]) & (!g181)) + ((!g25) & (!g120) & (g12) & (!sk[2]) & (g181)) + ((!g25) & (g120) & (g12) & (!sk[2]) & (!g181)));
	assign g241 = (((!g59) & (!sk[3]) & (g29) & (!g239) & (!g240)) + ((!g59) & (!sk[3]) & (!g29) & (g239) & (!g240)) + ((!g59) & (sk[3]) & (!g29) & (!g239) & (!g240)) + ((g59) & (!sk[3]) & (g29) & (!g239) & (!g240)));
	assign g242 = (((!g6) & (g88) & (!g238) & (!sk[4]) & (!g241)) + ((!g6) & (!g88) & (g238) & (!sk[4]) & (!g241)) + ((!g6) & (!g88) & (!g238) & (sk[4]) & (g241)) + ((!g6) & (!g88) & (!g238) & (sk[4]) & (g241)));
	assign g243 = (((!sk[5]) & (!g25) & (g36)) + ((sk[5]) & (!g25) & (!g36)));
	assign g244 = (((!g63) & (!sk[6]) & (!g51) & (g134)) + ((g63) & (!sk[6]) & (g51) & (g134)));
	assign g245 = (((!g2) & (g24) & (!sk[7]) & (!g32) & (!g244)) + ((!g2) & (!g24) & (!sk[7]) & (g32) & (!g244)) + ((!g2) & (g24) & (!sk[7]) & (!g32) & (!g244)) + ((!g2) & (!g24) & (sk[7]) & (!g32) & (!g244)) + ((!g2) & (!g24) & (!sk[7]) & (g32) & (!g244)));
	assign g246 = (((!i_6_) & (i_8_) & (!sk[8]) & (!g243) & (!g245)) + ((!i_6_) & (!i_8_) & (!sk[8]) & (g243) & (!g245)) + ((i_6_) & (!i_8_) & (sk[8]) & (!g243) & (g245)) + ((!i_6_) & (!i_8_) & (sk[8]) & (!g243) & (g245)) + ((!i_6_) & (!i_8_) & (sk[8]) & (!g243) & (g245)));
	assign g247 = (((g35) & (!sk[9]) & (!g42) & (!g25) & (!g23) & (!g3)) + ((!g35) & (!sk[9]) & (!g42) & (g25) & (!g23) & (!g3)) + ((!g35) & (!sk[9]) & (g42) & (!g25) & (g23) & (!g3)) + ((g35) & (!sk[9]) & (g42) & (!g25) & (!g23) & (g3)) + ((!g35) & (sk[9]) & (!g42) & (!g25) & (!g23) & (g3)));
	assign g248 = (((!g45) & (!g38) & (g29) & (!sk[10]) & (!g121)) + ((!g45) & (g38) & (!g29) & (!sk[10]) & (!g121)) + ((!g45) & (!g38) & (g29) & (!sk[10]) & (!g121)) + ((!g45) & (!g38) & (!g29) & (sk[10]) & (g121)));
	assign g249 = (((g21) & (!g8) & (!g25) & (!g247) & (!sk[11]) & (!g248)) + ((!g21) & (!g8) & (g25) & (!g247) & (!sk[11]) & (!g248)) + ((!g21) & (g8) & (!g25) & (g247) & (!sk[11]) & (!g248)) + ((g21) & (!g8) & (!g25) & (!g247) & (!sk[11]) & (!g248)) + ((!g21) & (!g8) & (g25) & (!g247) & (!sk[11]) & (!g248)) + ((!g21) & (!g8) & (!g25) & (!g247) & (sk[11]) & (!g248)));
	assign g250 = (((i_3_) & (!i_4_) & (!g27) & (!i_6_) & (!sk[12]) & (!i_8_)) + ((!i_3_) & (!i_4_) & (g27) & (!i_6_) & (!sk[12]) & (!i_8_)) + ((!i_3_) & (i_4_) & (!g27) & (i_6_) & (!sk[12]) & (!i_8_)) + ((i_3_) & (!i_4_) & (!g27) & (i_6_) & (!sk[12]) & (!i_8_)));
	assign g251 = (((i_3_) & (!sk[13]) & (!i_0_) & (!i_1_) & (!g219) & (!g250)) + ((!i_3_) & (!sk[13]) & (!i_0_) & (i_1_) & (!g219) & (!g250)) + ((i_3_) & (!sk[13]) & (!i_0_) & (!i_1_) & (!g219) & (!g250)) + ((!i_3_) & (!sk[13]) & (i_0_) & (!i_1_) & (g219) & (!g250)) + ((!i_3_) & (sk[13]) & (!i_0_) & (!i_1_) & (!g219) & (!g250)) + ((!i_3_) & (!sk[13]) & (i_0_) & (i_1_) & (!g219) & (!g250)) + ((!i_3_) & (!sk[13]) & (!i_0_) & (i_1_) & (!g219) & (!g250)));
	assign g252 = (((!g27) & (!g28) & (!sk[14]) & (g45)) + ((!g27) & (g28) & (sk[14]) & (!g45)));
	assign g253 = (((!sk[15]) & (g48) & (!g57) & (!g33) & (!g16) & (!g252)) + ((!sk[15]) & (!g48) & (!g57) & (g33) & (!g16) & (!g252)) + ((!sk[15]) & (!g48) & (g57) & (!g33) & (g16) & (!g252)) + ((sk[15]) & (!g48) & (!g57) & (!g33) & (!g16) & (!g252)) + ((sk[15]) & (!g48) & (!g57) & (!g33) & (!g16) & (!g252)) + ((sk[15]) & (!g48) & (!g57) & (!g33) & (!g16) & (!g252)) + ((sk[15]) & (!g48) & (!g57) & (!g33) & (!g16) & (!g252)));
	assign g254 = (((!sk[16]) & (g127) & (!g6) & (!g5) & (!g251) & (!g253)) + ((!sk[16]) & (!g127) & (!g6) & (g5) & (!g251) & (!g253)) + ((!sk[16]) & (!g127) & (g6) & (!g5) & (g251) & (!g253)) + ((sk[16]) & (!g127) & (!g6) & (!g5) & (g251) & (g253)) + ((sk[16]) & (!g127) & (!g6) & (!g5) & (g251) & (g253)) + ((sk[16]) & (!g127) & (!g6) & (!g5) & (g251) & (g253)));
	assign g255 = (((g14) & (!g1) & (!g12) & (!g3) & (!sk[17]) & (!g225)) + ((!g14) & (!g1) & (g12) & (!g3) & (!sk[17]) & (!g225)) + ((!g14) & (!g1) & (g12) & (g3) & (!sk[17]) & (!g225)) + ((!g14) & (g1) & (!g12) & (g3) & (!sk[17]) & (!g225)) + ((g14) & (!g1) & (!g12) & (!g3) & (!sk[17]) & (g225)));
	assign g256 = (((!g25) & (!sk[18]) & (!g120) & (g23)) + ((!g25) & (sk[18]) & (g120) & (!g23)));
	assign g257 = (((g8) & (!g1) & (!g22) & (!g105) & (!sk[19]) & (!g256)) + ((!g8) & (!g1) & (g22) & (!g105) & (!sk[19]) & (!g256)) + ((!g8) & (g1) & (!g22) & (g105) & (!sk[19]) & (!g256)) + ((!g8) & (g1) & (!g22) & (g105) & (!sk[19]) & (!g256)) + ((!g8) & (!g1) & (!g22) & (!g105) & (sk[19]) & (!g256)) + ((!g8) & (g1) & (!g22) & (!g105) & (sk[19]) & (!g256)) + ((!g8) & (!g1) & (!g22) & (g105) & (sk[19]) & (!g256)));
	assign g258 = (((g28) & (!g70) & (!g189) & (!g167) & (!sk[20]) & (!g230)) + ((!g28) & (!g70) & (g189) & (!g167) & (!sk[20]) & (!g230)) + ((!g28) & (!g70) & (!g189) & (!g167) & (sk[20]) & (!g230)) + ((!g28) & (g70) & (!g189) & (g167) & (!sk[20]) & (!g230)) + ((!g28) & (!g70) & (!g189) & (!g167) & (sk[20]) & (!g230)) + ((!g28) & (!g70) & (!g189) & (!g167) & (sk[20]) & (!g230)) + ((!g28) & (!g70) & (!g189) & (!g167) & (sk[20]) & (!g230)));
	assign g259 = (((!sk[21]) & (!g45) & (g6) & (!g110) & (!g141)) + ((!sk[21]) & (!g45) & (!g6) & (g110) & (!g141)) + ((!sk[21]) & (!g45) & (g6) & (g110) & (!g141)) + ((sk[21]) & (!g45) & (!g6) & (!g110) & (g141)));
	assign g260 = (((!sk[22]) & (g24) & (!g36) & (!g60) & (!g4) & (!g259)) + ((!sk[22]) & (!g24) & (!g36) & (g60) & (!g4) & (!g259)) + ((!sk[22]) & (g24) & (!g36) & (!g60) & (!g4) & (!g259)) + ((!sk[22]) & (!g24) & (g36) & (!g60) & (g4) & (!g259)) + ((sk[22]) & (!g24) & (!g36) & (!g60) & (!g4) & (!g259)) + ((!sk[22]) & (!g24) & (g36) & (g60) & (!g4) & (!g259)));
	assign g261 = (((g83) & (!g255) & (!sk[23]) & (!g257) & (!g258) & (!g260)) + ((!g83) & (!g255) & (!sk[23]) & (g257) & (!g258) & (!g260)) + ((!g83) & (g255) & (!sk[23]) & (!g257) & (g258) & (!g260)) + ((!g83) & (!g255) & (!sk[23]) & (g257) & (g258) & (g260)));
	assign g262 = (((g237) & (g242) & (g246) & (g249) & (g254) & (g261)));
	assign g263 = (((g157) & (g206) & (g211) & (g234) & (g236) & (g262)));
	assign g264 = (((!g11) & (g42) & (!g23) & (!g13) & (g60) & (!g38)) + ((!g11) & (!g42) & (!g23) & (!g13) & (!g60) & (!g38)));
	assign g265 = (((!sk[27]) & (!g27) & (!i_6_) & (g47)) + ((!sk[27]) & (!g27) & (!i_6_) & (g47)));
	assign g266 = (((!g11) & (g12) & (!sk[28]) & (!g71) & (!g265)) + ((!g11) & (g12) & (!sk[28]) & (g71) & (!g265)) + ((!g11) & (!g12) & (!sk[28]) & (g71) & (!g265)) + ((!g11) & (!g12) & (sk[28]) & (!g71) & (g265)));
	assign g267 = (((g27) & (!g35) & (!g36) & (!g110) & (!sk[29]) & (!g194)) + ((!g27) & (!g35) & (g36) & (!g110) & (!sk[29]) & (!g194)) + ((!g27) & (g35) & (!g36) & (g110) & (!sk[29]) & (!g194)) + ((!g27) & (!g35) & (!g36) & (!g110) & (sk[29]) & (g194)));
	assign g268 = (((!g24) & (!sk[30]) & (g225)) + ((!g24) & (!sk[30]) & (g225)));
	assign g269 = (((!i_7_) & (g28) & (g75) & (!sk[31]) & (!g268)) + ((!i_7_) & (g28) & (!g75) & (!sk[31]) & (!g268)) + ((!i_7_) & (!g28) & (g75) & (!sk[31]) & (!g268)) + ((i_7_) & (!g28) & (!g75) & (sk[31]) & (g268)));
	assign g270 = (((!sk[32]) & (!g1) & (g6) & (!g36) & (!g49)) + ((!sk[32]) & (!g1) & (!g6) & (g36) & (!g49)) + ((!sk[32]) & (!g1) & (g6) & (!g36) & (g49)) + ((!sk[32]) & (!g1) & (g6) & (!g36) & (!g49)));
	assign g271 = (((!g27) & (!g45) & (!g1) & (!g23) & (g4) & (!g189)) + ((!g27) & (!g45) & (!g1) & (!g23) & (!g4) & (g189)) + ((!g27) & (!g45) & (!g1) & (!g23) & (!g4) & (!g189)));
	assign g272 = (((!g48) & (g105) & (!g270) & (!sk[34]) & (!g271)) + ((!g48) & (!g105) & (g270) & (!sk[34]) & (!g271)) + ((!g48) & (g105) & (!g270) & (!sk[34]) & (!g271)) + ((!g48) & (!g105) & (!g270) & (sk[34]) & (!g271)));
	assign g273 = (((g8) & (!sk[35]) & (!g77) & (!g200) & (!g269) & (!g272)) + ((!g8) & (!sk[35]) & (!g77) & (g200) & (!g269) & (!g272)) + ((!g8) & (!sk[35]) & (g77) & (!g200) & (g269) & (!g272)) + ((!g8) & (sk[35]) & (!g77) & (!g200) & (!g269) & (g272)) + ((!g8) & (sk[35]) & (!g77) & (!g200) & (!g269) & (g272)));
	assign g274 = (((g264) & (!sk[36]) & (!g266) & (!g267) & (!g215) & (!g273)) + ((!g264) & (!sk[36]) & (!g266) & (g267) & (!g215) & (!g273)) + ((!g264) & (!sk[36]) & (g266) & (!g267) & (g215) & (!g273)) + ((!g264) & (sk[36]) & (!g266) & (!g267) & (g215) & (g273)));
	assign g275 = (((g27) & (!i_7_) & (!sk[37]) & (!i_8_) & (!g36) & (!g100)) + ((!g27) & (!i_7_) & (!sk[37]) & (i_8_) & (!g36) & (!g100)) + ((!g27) & (i_7_) & (!sk[37]) & (!i_8_) & (g36) & (!g100)) + ((!g27) & (i_7_) & (!sk[37]) & (i_8_) & (!g36) & (g100)) + ((!g27) & (i_7_) & (sk[37]) & (!i_8_) & (!g36) & (!g100)));
	assign g276 = (((!sk[38]) & (g28) & (!g42) & (!g23) & (!g3) & (!g91)) + ((!sk[38]) & (!g28) & (!g42) & (g23) & (!g3) & (!g91)) + ((!sk[38]) & (!g28) & (g42) & (!g23) & (g3) & (!g91)) + ((!sk[38]) & (g28) & (g42) & (!g23) & (g3) & (!g91)) + ((sk[38]) & (!g28) & (!g42) & (!g23) & (!g3) & (g91)));
	assign g277 = (((g11) & (!g8) & (!g12) & (!sk[39]) & (!g13) & (!g184)) + ((!g11) & (!g8) & (g12) & (!sk[39]) & (!g13) & (!g184)) + ((!g11) & (g8) & (!g12) & (!sk[39]) & (g13) & (!g184)) + ((!g11) & (!g8) & (g12) & (!sk[39]) & (!g13) & (!g184)) + ((!g11) & (g8) & (!g12) & (sk[39]) & (!g13) & (g184)));
	assign g278 = (((!sk[40]) & (!g35) & (!g46) & (g158)) + ((!sk[40]) & (g35) & (!g46) & (g158)) + ((sk[40]) & (g35) & (g46) & (!g158)));
	assign g279 = (((!g38) & (g94) & (!sk[41]) & (!g265) & (!g167)) + ((!g38) & (!g94) & (!sk[41]) & (g265) & (!g167)) + ((!g38) & (!g94) & (!sk[41]) & (g265) & (!g167)) + ((!g38) & (g94) & (!sk[41]) & (!g265) & (g167)));
	assign g280 = (((g25) & (!sk[42]) & (!g6) & (!g32) & (!g121) & (!g252)) + ((!g25) & (!sk[42]) & (!g6) & (g32) & (!g121) & (!g252)) + ((!g25) & (!sk[42]) & (g6) & (!g32) & (g121) & (!g252)) + ((!g25) & (sk[42]) & (!g6) & (!g32) & (!g121) & (!g252)) + ((g25) & (!sk[42]) & (!g6) & (!g32) & (!g121) & (!g252)) + ((!g25) & (!sk[42]) & (!g6) & (g32) & (!g121) & (!g252)));
	assign g281 = (((!sk[43]) & (!g35) & (g6) & (!g117) & (!g161)) + ((!sk[43]) & (!g35) & (!g6) & (g117) & (!g161)) + ((!sk[43]) & (g35) & (!g6) & (g117) & (!g161)) + ((!sk[43]) & (!g35) & (g6) & (!g117) & (g161)));
	assign g282 = (((g277) & (!sk[44]) & (!g278) & (!g279) & (!g280) & (!g281)) + ((!g277) & (!sk[44]) & (!g278) & (g279) & (!g280) & (!g281)) + ((!g277) & (!sk[44]) & (g278) & (!g279) & (g280) & (!g281)) + ((!g277) & (sk[44]) & (!g278) & (!g279) & (g280) & (!g281)));
	assign g283 = (((i_0_) & (!g135) & (!g275) & (!g276) & (!sk[45]) & (!g282)) + ((!i_0_) & (!g135) & (g275) & (!g276) & (!sk[45]) & (!g282)) + ((!i_0_) & (g135) & (!g275) & (g276) & (!sk[45]) & (!g282)) + ((!i_0_) & (!g135) & (!g275) & (!g276) & (sk[45]) & (g282)) + ((!i_0_) & (!g135) & (!g275) & (!g276) & (sk[45]) & (g282)));
	assign g284 = (((!sk[46]) & (!g27) & (!g137) & (g15)) + ((!sk[46]) & (!g27) & (g137) & (g15)));
	assign g285 = (((!i_6_) & (i_8_) & (!g1) & (!sk[47]) & (!g32)) + ((!i_6_) & (!i_8_) & (g1) & (!sk[47]) & (!g32)) + ((!i_6_) & (!i_8_) & (!g1) & (sk[47]) & (g32)));
	assign g286 = (((!g2) & (!g26) & (!sk[48]) & (g155)) + ((!g2) & (!g26) & (sk[48]) & (!g155)) + ((!g2) & (!g26) & (sk[48]) & (!g155)));
	assign g287 = (((g25) & (!g194) & (!g212) & (!g285) & (!sk[49]) & (!g286)) + ((!g25) & (!g194) & (g212) & (!g285) & (!sk[49]) & (!g286)) + ((!g25) & (g194) & (!g212) & (g285) & (!sk[49]) & (!g286)) + ((g25) & (!g194) & (!g212) & (!g285) & (!sk[49]) & (g286)) + ((!g25) & (!g194) & (!g212) & (!g285) & (sk[49]) & (g286)));
	assign g288 = (((!g28) & (g12) & (g184) & (!sk[50]) & (!g243)) + ((!g28) & (g12) & (!g184) & (!sk[50]) & (!g243)) + ((!g28) & (!g12) & (g184) & (!sk[50]) & (!g243)) + ((g28) & (!g12) & (!g184) & (sk[50]) & (g243)));
	assign g289 = (((g13) & (!g123) & (!sk[51]) & (!g284) & (!g287) & (!g288)) + ((!g13) & (!g123) & (!sk[51]) & (g284) & (!g287) & (!g288)) + ((!g13) & (g123) & (!sk[51]) & (!g284) & (g287) & (!g288)) + ((g13) & (!g123) & (!sk[51]) & (!g284) & (g287) & (!g288)) + ((!g13) & (!g123) & (sk[51]) & (!g284) & (g287) & (!g288)));
	assign g290 = (((!g42) & (!sk[52]) & (!g2) & (g38)) + ((g42) & (sk[52]) & (g2) & (!g38)));
	assign g291 = (((!g48) & (g181) & (!sk[53]) & (!g244) & (!g290)) + ((!g48) & (!g181) & (!sk[53]) & (g244) & (!g290)) + ((!g48) & (!g181) & (sk[53]) & (!g244) & (!g290)) + ((!g48) & (!g181) & (sk[53]) & (!g244) & (!g290)));
	assign g292 = (((!g27) & (!sk[54]) & (i_6_) & (!i_8_) & (!g21)) + ((!g27) & (!sk[54]) & (!i_6_) & (i_8_) & (!g21)) + ((!g27) & (!sk[54]) & (i_6_) & (!i_8_) & (!g21)));
	assign g293 = (((!sk[55]) & (g27) & (!g35) & (!g45) & (!g6) & (!g84)) + ((!sk[55]) & (!g27) & (!g35) & (g45) & (!g6) & (!g84)) + ((sk[55]) & (!g27) & (g35) & (!g45) & (!g6) & (g84)) + ((sk[55]) & (!g27) & (!g35) & (!g45) & (g6) & (!g84)) + ((!sk[55]) & (!g27) & (g35) & (!g45) & (g6) & (!g84)));
	assign g294 = (((!sk[56]) & (!g28) & (!g45) & (g24)) + ((sk[56]) & (g28) & (!g45) & (!g24)));
	assign g295 = (((!i_5_) & (!g35) & (!g42) & (!g5) & (!g121) & (!g294)) + ((!i_5_) & (!g35) & (!g42) & (!g5) & (!g121) & (!g294)) + ((!i_5_) & (!g35) & (!g42) & (!g5) & (!g121) & (!g294)) + ((i_5_) & (!g35) & (!g42) & (!g5) & (!g121) & (!g294)));
	assign g296 = (((!sk[58]) & (!g8) & (g243)) + ((!sk[58]) & (g8) & (g243)));
	assign g297 = (((!sk[59]) & (i_3_) & (!i_5_) & (!g35) & (!g14) & (!g85)) + ((!sk[59]) & (!i_3_) & (!i_5_) & (g35) & (!g14) & (!g85)) + ((!sk[59]) & (!i_3_) & (!i_5_) & (g35) & (!g14) & (!g85)) + ((!sk[59]) & (!i_3_) & (i_5_) & (!g35) & (g14) & (!g85)) + ((sk[59]) & (!i_3_) & (!i_5_) & (!g35) & (g14) & (g85)));
	assign g298 = (((g23) & (!g24) & (!g70) & (!g296) & (!sk[60]) & (!g297)) + ((!g23) & (!g24) & (g70) & (!g296) & (!sk[60]) & (!g297)) + ((g23) & (g24) & (!g70) & (!g296) & (!sk[60]) & (!g297)) + ((!g23) & (g24) & (!g70) & (g296) & (!sk[60]) & (!g297)) + ((g23) & (!g24) & (!g70) & (!g296) & (!sk[60]) & (!g297)) + ((!g23) & (g24) & (!g70) & (!g296) & (sk[60]) & (!g297)) + ((!g23) & (!g24) & (!g70) & (!g296) & (sk[60]) & (!g297)));
	assign g299 = (((!g292) & (!sk[61]) & (g293) & (!g295) & (!g298)) + ((!g292) & (!sk[61]) & (!g293) & (g295) & (!g298)) + ((!g292) & (!sk[61]) & (!g293) & (g295) & (g298)));
	assign g300 = (((g164) & (!sk[62]) & (!g283) & (!g289) & (!g291) & (!g299)) + ((!g164) & (!sk[62]) & (!g283) & (g289) & (!g291) & (!g299)) + ((!g164) & (!sk[62]) & (g283) & (!g289) & (g291) & (!g299)) + ((g164) & (!sk[62]) & (g283) & (g289) & (g291) & (g299)));
	assign g301 = (((!sk[63]) & (i_6_) & (!g137) & (!g77) & (!g13) & (!g64)) + ((!sk[63]) & (!i_6_) & (!g137) & (g77) & (!g13) & (!g64)) + ((!sk[63]) & (!i_6_) & (g137) & (g77) & (!g13) & (!g64)) + ((!sk[63]) & (!i_6_) & (g137) & (!g77) & (g13) & (!g64)) + ((sk[63]) & (!i_6_) & (g137) & (!g77) & (!g13) & (g64)));
	assign g302 = (((i_6_) & (!sk[64]) & (!g21) & (!g1) & (!g137) & (!g59)) + ((!i_6_) & (!sk[64]) & (!g21) & (g1) & (!g137) & (!g59)) + ((!i_6_) & (!sk[64]) & (g21) & (!g1) & (g137) & (!g59)) + ((i_6_) & (!sk[64]) & (!g21) & (!g1) & (g137) & (!g59)) + ((!i_6_) & (sk[64]) & (!g21) & (!g1) & (g137) & (!g59)));
	assign g303 = (((!g27) & (!sk[65]) & (g63) & (!g38) & (!g96)) + ((!g27) & (!sk[65]) & (!g63) & (g38) & (!g96)) + ((!g27) & (!sk[65]) & (!g63) & (g38) & (!g96)) + ((!g27) & (sk[65]) & (!g63) & (!g38) & (!g96)) + ((g27) & (!sk[65]) & (g63) & (!g38) & (!g96)));
	assign g304 = (((g35) & (!g45) & (!g13) & (!sk[66]) & (!g4) & (!g243)) + ((!g35) & (!g45) & (g13) & (!sk[66]) & (!g4) & (!g243)) + ((g35) & (!g45) & (!g13) & (!sk[66]) & (!g4) & (g243)) + ((g35) & (!g45) & (!g13) & (!sk[66]) & (!g4) & (!g243)) + ((!g35) & (!g45) & (!g13) & (sk[66]) & (g4) & (!g243)) + ((!g35) & (g45) & (!g13) & (!sk[66]) & (g4) & (!g243)));
	assign g305 = (((!g2) & (g6) & (!sk[67]) & (!g75) & (!g71)) + ((g2) & (!g6) & (!sk[67]) & (g75) & (!g71)) + ((!g2) & (!g6) & (!sk[67]) & (g75) & (!g71)) + ((!g2) & (g6) & (!sk[67]) & (!g75) & (g71)));
	assign g306 = (((g23) & (!g184) & (!sk[68]) & (!g304) & (!g607) & (!g305)) + ((!g23) & (!g184) & (!sk[68]) & (g304) & (!g607) & (!g305)) + ((!g23) & (g184) & (!sk[68]) & (!g304) & (g607) & (!g305)) + ((g23) & (!g184) & (!sk[68]) & (!g304) & (g607) & (!g305)) + ((!g23) & (!g184) & (sk[68]) & (!g304) & (g607) & (!g305)));
	assign g307 = (((g11) & (!sk[69]) & (!g67) & (!g302) & (!g303) & (!g306)) + ((!g11) & (!sk[69]) & (!g67) & (g302) & (!g303) & (!g306)) + ((!g11) & (!sk[69]) & (g67) & (!g302) & (g303) & (!g306)) + ((g11) & (!sk[69]) & (!g67) & (!g302) & (g303) & (g306)) + ((!g11) & (sk[69]) & (!g67) & (!g302) & (g303) & (g306)));
	assign g308 = (((!i_3_) & (!i_4_) & (!i_0_) & (i_2_) & (!g12) & (g219)) + ((i_3_) & (!i_4_) & (!i_0_) & (i_2_) & (g12) & (!g219)));
	assign g309 = (((!g42) & (g23) & (!sk[71]) & (!g194) & (!g98)) + ((g42) & (!g23) & (!sk[71]) & (g194) & (!g98)) + ((!g42) & (!g23) & (!sk[71]) & (g194) & (!g98)) + ((!g42) & (!g23) & (sk[71]) & (!g194) & (g98)));
	assign g310 = (((!i_6_) & (i_7_) & (!sk[72]) & (!g129) & (!g309)) + ((!i_6_) & (!i_7_) & (!sk[72]) & (g129) & (!g309)) + ((!i_6_) & (i_7_) & (!sk[72]) & (!g129) & (!g309)) + ((!i_6_) & (!i_7_) & (sk[72]) & (!g129) & (!g309)) + ((!i_6_) & (!i_7_) & (!sk[72]) & (g129) & (!g309)));
	assign g311 = (((g2) & (!sk[73]) & (!g23) & (!g59) & (!g13) & (!g84)) + ((!g2) & (!sk[73]) & (!g23) & (g59) & (!g13) & (!g84)) + ((!g2) & (!sk[73]) & (g23) & (!g59) & (g13) & (!g84)) + ((g2) & (!sk[73]) & (!g23) & (!g59) & (!g13) & (!g84)) + ((!g2) & (sk[73]) & (!g23) & (!g59) & (!g13) & (g84)));
	assign g312 = (((i_3_) & (!sk[74]) & (!i_4_) & (!g28) & (!g24) & (!g311)) + ((!i_3_) & (!sk[74]) & (!i_4_) & (g28) & (!g24) & (!g311)) + ((!i_3_) & (!sk[74]) & (i_4_) & (!g28) & (g24) & (!g311)) + ((!i_3_) & (sk[74]) & (!i_4_) & (!g28) & (!g24) & (!g311)) + ((!i_3_) & (sk[74]) & (i_4_) & (!g28) & (!g24) & (!g311)) + ((!i_3_) & (sk[74]) & (!i_4_) & (!g28) & (!g24) & (!g311)) + ((!i_3_) & (!sk[74]) & (!i_4_) & (g28) & (g24) & (!g311)));
	assign g313 = (((g25) & (!sk[75]) & (!g12) & (!g32) & (!g9) & (!g116)) + ((!g25) & (!sk[75]) & (!g12) & (g32) & (!g9) & (!g116)) + ((!g25) & (!sk[75]) & (g12) & (g32) & (!g9) & (!g116)) + ((!g25) & (!sk[75]) & (g12) & (!g32) & (g9) & (!g116)) + ((!g25) & (sk[75]) & (!g12) & (!g32) & (g9) & (g116)));
	assign g314 = (((g11) & (!g48) & (!g24) & (!g32) & (!sk[76]) & (!g9)) + ((!g11) & (!g48) & (g24) & (!g32) & (!sk[76]) & (!g9)) + ((!g11) & (g48) & (!g24) & (g32) & (!sk[76]) & (!g9)) + ((!g11) & (!g48) & (!g24) & (!g32) & (sk[76]) & (g9)));
	assign g315 = (((!g1) & (!sk[77]) & (!g32) & (g37)) + ((!g1) & (!sk[77]) & (g32) & (g37)));
	assign g316 = (((!g6) & (!sk[78]) & (!g105) & (g315)) + ((!g6) & (sk[78]) & (!g105) & (!g315)) + ((!g6) & (sk[78]) & (g105) & (!g315)));
	assign g317 = (((g48) & (!sk[79]) & (!g313) & (!g314) & (!g52) & (!g316)) + ((!g48) & (!sk[79]) & (!g313) & (g314) & (!g52) & (!g316)) + ((!g48) & (!sk[79]) & (g313) & (!g314) & (g52) & (!g316)) + ((!g48) & (sk[79]) & (!g313) & (!g314) & (!g52) & (g316)) + ((!g48) & (sk[79]) & (!g313) & (!g314) & (!g52) & (g316)));
	assign g318 = (((!g168) & (g310) & (!sk[80]) & (!g312) & (!g317)) + ((!g168) & (!g310) & (!sk[80]) & (g312) & (!g317)) + ((!g168) & (g310) & (!sk[80]) & (g312) & (g317)));
	assign g319 = (((!sk[81]) & (g301) & (!g211) & (!g307) & (!g308) & (!g318)) + ((!sk[81]) & (!g301) & (!g211) & (g307) & (!g308) & (!g318)) + ((!sk[81]) & (!g301) & (g211) & (!g307) & (g308) & (!g318)) + ((!sk[81]) & (!g301) & (g211) & (g307) & (!g308) & (g318)));
	assign g320 = (((g90) & (g224) & (g274) & (g618) & (g300) & (g319)));
	assign g321 = (((!i_6_) & (i_7_) & (!i_8_) & (!g26) & (g243) & (!g268)) + ((!i_6_) & (i_7_) & (i_8_) & (!g26) & (!g243) & (g268)) + ((i_6_) & (!i_7_) & (!i_8_) & (g26) & (!g243) & (!g268)));
	assign g322 = (((g27) & (!g45) & (!g1) & (!g6) & (!sk[84]) & (!g16)) + ((!g27) & (!g45) & (g1) & (!g6) & (!sk[84]) & (!g16)) + ((!g27) & (g45) & (!g1) & (g6) & (!sk[84]) & (!g16)) + ((!g27) & (!g45) & (!g1) & (!g6) & (sk[84]) & (g16)) + ((!g27) & (!g45) & (!g1) & (g6) & (sk[84]) & (!g16)));
	assign g323 = (((!sk[85]) & (g264) & (!g279) & (!g596) & (!g321) & (!g322)) + ((!sk[85]) & (!g264) & (!g279) & (g596) & (!g321) & (!g322)) + ((!sk[85]) & (!g264) & (g279) & (!g596) & (g321) & (!g322)) + ((!sk[85]) & (!g264) & (!g279) & (g596) & (!g321) & (!g322)));
	assign g324 = (((g28) & (!g48) & (g189) & (!sk[86]) & (!g184)) + ((!g28) & (g48) & (!g189) & (!sk[86]) & (!g184)) + ((!g28) & (!g48) & (g189) & (!sk[86]) & (!g184)) + ((!g28) & (g48) & (!g189) & (!sk[86]) & (g184)));
	assign g325 = (((!g137) & (!sk[87]) & (!g134) & (g230)) + ((g137) & (!sk[87]) & (g134) & (g230)));
	assign g326 = (((g35) & (!g25) & (!g59) & (!g4) & (!sk[88]) & (!g325)) + ((!g35) & (!g25) & (g59) & (!g4) & (!sk[88]) & (!g325)) + ((!g35) & (g25) & (!g59) & (g4) & (!sk[88]) & (!g325)) + ((!g35) & (!g25) & (g59) & (!g4) & (!sk[88]) & (!g325)) + ((!g35) & (!g25) & (!g59) & (!g4) & (sk[88]) & (!g325)) + ((!g35) & (g25) & (!g59) & (!g4) & (sk[88]) & (!g325)));
	assign g327 = (((g35) & (!sk[89]) & (!g181) & (!g276) & (!g324) & (!g326)) + ((!g35) & (!sk[89]) & (!g181) & (g276) & (!g324) & (!g326)) + ((!g35) & (!sk[89]) & (g181) & (!g276) & (g324) & (!g326)) + ((!g35) & (sk[89]) & (!g181) & (!g276) & (!g324) & (g326)) + ((!g35) & (sk[89]) & (!g181) & (!g276) & (!g324) & (g326)));
	assign g328 = (((!i_6_) & (!sk[90]) & (g14) & (!g26) & (!g99)) + ((!i_6_) & (!sk[90]) & (!g14) & (g26) & (!g99)) + ((!i_6_) & (!sk[90]) & (g14) & (g26) & (!g99)) + ((i_6_) & (!sk[90]) & (g14) & (!g26) & (g99)));
	assign g329 = (((g45) & (!sk[91]) & (!g6) & (!g24) & (!g67) & (!g91)) + ((!g45) & (!sk[91]) & (!g6) & (g24) & (!g67) & (!g91)) + ((!g45) & (sk[91]) & (!g6) & (!g24) & (g67) & (!g91)) + ((!g45) & (sk[91]) & (g6) & (!g24) & (!g67) & (!g91)) + ((!g45) & (!sk[91]) & (g6) & (!g24) & (g67) & (!g91)) + ((!g45) & (sk[91]) & (g6) & (!g24) & (!g67) & (g91)));
	assign g330 = (((g32) & (!g29) & (!g193) & (!g328) & (!sk[92]) & (!g329)) + ((!g32) & (!g29) & (g193) & (!g328) & (!sk[92]) & (!g329)) + ((!g32) & (g29) & (!g193) & (g328) & (!sk[92]) & (!g329)) + ((!g32) & (!g29) & (!g193) & (!g328) & (sk[92]) & (!g329)) + ((!g32) & (!g29) & (!g193) & (!g328) & (sk[92]) & (!g329)));
	assign g331 = (((!g14) & (!g64) & (!sk[93]) & (g230)) + ((g14) & (g64) & (!sk[93]) & (g230)));
	assign g332 = (((!sk[94]) & (g45) & (!g2) & (!g49) & (!g7) & (!g331)) + ((!sk[94]) & (!g45) & (!g2) & (g49) & (!g7) & (!g331)) + ((!sk[94]) & (!g45) & (g2) & (!g49) & (g7) & (!g331)) + ((!sk[94]) & (g45) & (!g2) & (!g49) & (!g7) & (!g331)) + ((!sk[94]) & (g45) & (!g2) & (!g49) & (!g7) & (!g331)) + ((sk[94]) & (!g45) & (!g2) & (!g49) & (!g7) & (!g331)) + ((!sk[94]) & (!g45) & (!g2) & (g49) & (!g7) & (!g331)));
	assign g333 = (((i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (i_8_)) + ((i_3_) & (i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (!i_8_)));
	assign g334 = (((!i_3_) & (g27) & (!i_6_) & (!sk[96]) & (!g333)) + ((!i_3_) & (!g27) & (i_6_) & (!sk[96]) & (!g333)) + ((i_3_) & (!g27) & (!i_6_) & (sk[96]) & (g333)));
	assign g335 = (((!g11) & (!g35) & (!g28) & (g25) & (!g38) & (!g334)) + ((g11) & (!g35) & (!g28) & (!g25) & (!g38) & (!g334)) + ((!g11) & (!g35) & (!g28) & (!g25) & (!g38) & (!g334)) + ((g11) & (!g35) & (!g28) & (!g25) & (g38) & (!g334)) + ((!g11) & (!g35) & (!g28) & (!g25) & (g38) & (!g334)));
	assign g336 = (((i_3_) & (!sk[98]) & (!g21) & (!g42) & (!g8) & (!g7)) + ((!i_3_) & (!sk[98]) & (!g21) & (g42) & (!g8) & (!g7)) + ((!i_3_) & (!sk[98]) & (g21) & (!g42) & (g8) & (!g7)) + ((i_3_) & (!sk[98]) & (!g21) & (g42) & (g8) & (!g7)) + ((!i_3_) & (sk[98]) & (!g21) & (!g42) & (!g8) & (g7)));
	assign g337 = (((!sk[99]) & (i_6_) & (!i_7_) & (!i_8_) & (!g70) & (!g184)) + ((!sk[99]) & (!i_6_) & (!i_7_) & (i_8_) & (!g70) & (!g184)) + ((!sk[99]) & (!i_6_) & (i_7_) & (!i_8_) & (g70) & (!g184)) + ((!sk[99]) & (i_6_) & (!i_7_) & (!i_8_) & (g70) & (!g184)) + ((sk[99]) & (!i_6_) & (i_7_) & (!i_8_) & (!g70) & (g184)));
	assign g338 = (((!sk[100]) & (!g46) & (!g48) & (g60)) + ((!sk[100]) & (g46) & (!g48) & (g60)) + ((sk[100]) & (g46) & (g48) & (!g60)));
	assign g339 = (((g2) & (!g98) & (!g252) & (!g337) & (!sk[101]) & (!g338)) + ((!g2) & (!g98) & (g252) & (!g337) & (!sk[101]) & (!g338)) + ((!g2) & (g98) & (!g252) & (g337) & (!sk[101]) & (!g338)) + ((!g2) & (!g98) & (!g252) & (!g337) & (sk[101]) & (!g338)) + ((!g2) & (!g98) & (!g252) & (!g337) & (sk[101]) & (!g338)));
	assign g340 = (((g312) & (!g332) & (!sk[102]) & (!g335) & (!g336) & (!g339)) + ((!g312) & (!g332) & (!sk[102]) & (g335) & (!g336) & (!g339)) + ((!g312) & (g332) & (!sk[102]) & (!g335) & (g336) & (!g339)) + ((g312) & (g332) & (!sk[102]) & (g335) & (!g336) & (g339)));
	assign g341 = (((!sk[103]) & (g119) & (!g206) & (!g327) & (!g330) & (!g340)) + ((!sk[103]) & (!g119) & (!g206) & (g327) & (!g330) & (!g340)) + ((!sk[103]) & (!g119) & (g206) & (!g327) & (g330) & (!g340)) + ((!sk[103]) & (g119) & (g206) & (g327) & (g330) & (g340)));
	assign g342 = (((i_0_) & (!g27) & (!g14) & (g135) & (!sk[104]) & (!g217)) + ((i_0_) & (!g27) & (!g14) & (!g135) & (!sk[104]) & (!g217)) + ((!i_0_) & (!g27) & (g14) & (!g135) & (!sk[104]) & (!g217)) + ((!i_0_) & (g27) & (!g14) & (g135) & (!sk[104]) & (!g217)) + ((!i_0_) & (!g27) & (g14) & (!g135) & (!sk[104]) & (g217)));
	assign g343 = (((!g27) & (g23) & (!g36) & (!sk[105]) & (!g285)) + ((!g27) & (!g23) & (g36) & (!sk[105]) & (!g285)) + ((!g27) & (g23) & (!g36) & (!sk[105]) & (!g285)) + ((!g27) & (!g23) & (g36) & (!sk[105]) & (!g285)) + ((g27) & (!g23) & (!g36) & (sk[105]) & (!g285)));
	assign g344 = (((!sk[106]) & (g21) & (!g6) & (!g23) & (!g24) & (!g129)) + ((!sk[106]) & (!g21) & (!g6) & (g23) & (!g24) & (!g129)) + ((!sk[106]) & (!g21) & (g6) & (!g23) & (g24) & (!g129)) + ((sk[106]) & (!g21) & (!g6) & (!g23) & (!g24) & (!g129)) + ((sk[106]) & (!g21) & (g6) & (!g23) & (!g24) & (g129)));
	assign g345 = (((i_5_) & (!i_6_) & (!i_7_) & (!i_8_) & (!sk[107]) & (!g5)) + ((!i_5_) & (!i_6_) & (i_7_) & (!i_8_) & (!sk[107]) & (!g5)) + ((!i_5_) & (i_6_) & (!i_7_) & (i_8_) & (!sk[107]) & (!g5)) + ((i_5_) & (!i_6_) & (i_7_) & (!i_8_) & (!sk[107]) & (g5)) + ((!i_5_) & (i_6_) & (!i_7_) & (!i_8_) & (sk[107]) & (g5)));
	assign g346 = (((!g28) & (!g42) & (!g38) & (g110) & (g159) & (!g345)) + ((!g28) & (g42) & (!g38) & (!g110) & (!g159) & (g345)) + ((g28) & (!g42) & (!g38) & (g110) & (!g159) & (!g345)));
	assign g347 = (((i_6_) & (!i_7_) & (!i_8_) & (g46) & (!g77) & (!g189)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g46) & (!g77) & (!g189)) + ((i_6_) & (!i_7_) & (i_8_) & (!g46) & (g77) & (!g189)) + ((i_6_) & (!i_7_) & (i_8_) & (!g46) & (!g77) & (g189)));
	assign g348 = (((!i_3_) & (i_4_) & (!sk[110]) & (!i_0_) & (!i_1_)) + ((!i_3_) & (!i_4_) & (!sk[110]) & (i_0_) & (!i_1_)) + ((i_3_) & (!i_4_) & (!sk[110]) & (i_0_) & (!i_1_)));
	assign g349 = (((!sk[111]) & (!g2) & (g161) & (!g296) & (!g348)) + ((!sk[111]) & (!g2) & (!g161) & (g296) & (!g348)) + ((sk[111]) & (!g2) & (!g161) & (!g296) & (!g348)) + ((sk[111]) & (!g2) & (!g161) & (!g296) & (!g348)));
	assign g350 = (((!sk[112]) & (g343) & (!g344) & (!g346) & (!g347) & (!g349)) + ((!sk[112]) & (!g343) & (!g344) & (g346) & (!g347) & (!g349)) + ((!sk[112]) & (!g343) & (g344) & (!g346) & (g347) & (!g349)) + ((!sk[112]) & (g343) & (!g344) & (!g346) & (!g347) & (g349)));
	assign g351 = (((!i_5_) & (!sk[113]) & (i_2_) & (!g48) & (!g219)) + ((!i_5_) & (!sk[113]) & (!i_2_) & (g48) & (!g219)) + ((!i_5_) & (!sk[113]) & (i_2_) & (!g48) & (!g219)) + ((!i_5_) & (sk[113]) & (!i_2_) & (!g48) & (!g219)) + ((i_5_) & (!sk[113]) & (!i_2_) & (g48) & (!g219)));
	assign g352 = (((!i_3_) & (!sk[114]) & (i_0_) & (!i_1_) & (!g351)) + ((!i_3_) & (!sk[114]) & (!i_0_) & (i_1_) & (!g351)) + ((!i_3_) & (!sk[114]) & (!i_0_) & (i_1_) & (!g351)));
	assign g353 = (((!g50) & (!sk[115]) & (i_6_) & (!i_7_) & (!g86)) + ((!g50) & (!sk[115]) & (!i_6_) & (i_7_) & (!g86)) + ((g50) & (!sk[115]) & (i_6_) & (!i_7_) & (g86)));
	assign g354 = (((g13) & (!g4) & (!g352) & (!sk[116]) & (!g125) & (!g353)) + ((!g13) & (!g4) & (g352) & (!sk[116]) & (!g125) & (!g353)) + ((!g13) & (g4) & (!g352) & (!sk[116]) & (g125) & (!g353)) + ((g13) & (!g4) & (!g352) & (!sk[116]) & (g125) & (!g353)) + ((!g13) & (!g4) & (!g352) & (sk[116]) & (g125) & (!g353)));
	assign g355 = (((g301) & (!g20) & (!g342) & (!sk[117]) & (!g350) & (!g354)) + ((!g301) & (!g20) & (g342) & (!sk[117]) & (!g350) & (!g354)) + ((!g301) & (g20) & (!g342) & (!sk[117]) & (g350) & (!g354)) + ((!g301) & (g20) & (!g342) & (!sk[117]) & (g350) & (g354)));
	assign g356 = (((g178) & (!g234) & (!sk[118]) & (!g323) & (!g341) & (!g355)) + ((!g178) & (!g234) & (!sk[118]) & (g323) & (!g341) & (!g355)) + ((!g178) & (g234) & (!sk[118]) & (!g323) & (g341) & (!g355)) + ((g178) & (g234) & (!sk[118]) & (g323) & (g341) & (g355)));
	assign g357 = (((!g6) & (g4) & (g110) & (!sk[119]) & (!g243)) + ((!g6) & (g4) & (!g110) & (!sk[119]) & (!g243)) + ((!g6) & (!g4) & (g110) & (!sk[119]) & (!g243)) + ((g6) & (!g4) & (!g110) & (sk[119]) & (g243)));
	assign g358 = (((!i_6_) & (i_7_) & (!g75) & (!sk[120]) & (!g357)) + ((!i_6_) & (!i_7_) & (g75) & (!sk[120]) & (!g357)) + ((!i_6_) & (i_7_) & (!g75) & (!sk[120]) & (!g357)) + ((!i_6_) & (!i_7_) & (!g75) & (sk[120]) & (!g357)) + ((!i_6_) & (!i_7_) & (!g75) & (sk[120]) & (!g357)));
	assign g359 = (((!sk[121]) & (!g21) & (g110)) + ((!sk[121]) & (!g21) & (g110)));
	assign g360 = (((!i_6_) & (!i_7_) & (i_8_) & (g73) & (!g184) & (!g359)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g73) & (g184) & (!g359)) + ((!i_6_) & (!i_7_) & (!i_8_) & (!g73) & (!g184) & (g359)));
	assign g361 = (((!sk[123]) & (g127) & (!i_2_) & (!i_6_) & (!g137) & (!g5)) + ((!sk[123]) & (!g127) & (!i_2_) & (i_6_) & (!g137) & (!g5)) + ((!sk[123]) & (!g127) & (i_2_) & (!i_6_) & (g137) & (!g5)) + ((!sk[123]) & (g127) & (i_2_) & (i_6_) & (g137) & (g5)) + ((!sk[123]) & (g127) & (!i_2_) & (!i_6_) & (g137) & (g5)));
	assign g362 = (((!sk[124]) & (g11) & (!g42) & (!g22) & (!g121) & (!g361)) + ((!sk[124]) & (!g11) & (!g42) & (g22) & (!g121) & (!g361)) + ((!sk[124]) & (!g11) & (g42) & (!g22) & (g121) & (!g361)) + ((!sk[124]) & (g11) & (!g42) & (!g22) & (!g121) & (!g361)) + ((!sk[124]) & (g11) & (!g42) & (!g22) & (!g121) & (!g361)) + ((sk[124]) & (!g11) & (!g42) & (!g22) & (!g121) & (!g361)) + ((!sk[124]) & (!g11) & (!g42) & (g22) & (!g121) & (!g361)));
	assign g363 = (((!i_4_) & (!sk[125]) & (i_5_) & (!g23) & (!g110)) + ((!i_4_) & (!sk[125]) & (!i_5_) & (g23) & (!g110)) + ((i_4_) & (!sk[125]) & (i_5_) & (!g23) & (g110)));
	assign g364 = (((!g21) & (!g6) & (!sk[126]) & (g24)) + ((!g21) & (g6) & (sk[126]) & (!g24)));
	assign g365 = (((g21) & (!sk[127]) & (!g38) & (!g7) & (!g265) & (!g364)) + ((!g21) & (!sk[127]) & (!g38) & (g7) & (!g265) & (!g364)) + ((!g21) & (!sk[127]) & (g38) & (!g7) & (g265) & (!g364)) + ((g21) & (!sk[127]) & (g38) & (!g7) & (!g265) & (!g364)) + ((g21) & (!sk[127]) & (!g38) & (!g7) & (!g265) & (!g364)) + ((!g21) & (sk[127]) & (!g38) & (!g7) & (!g265) & (!g364)) + ((!g21) & (!sk[127]) & (g38) & (g7) & (!g265) & (!g364)));
	assign g366 = (((!sk[0]) & (!g175) & (g256) & (!g363) & (!g365)) + ((!sk[0]) & (!g175) & (!g256) & (g363) & (!g365)) + ((sk[0]) & (!g175) & (!g256) & (!g363) & (g365)));
	assign g367 = (((!sk[1]) & (g202) & (!g358) & (!g360) & (!g362) & (!g366)) + ((!sk[1]) & (!g202) & (!g358) & (g360) & (!g362) & (!g366)) + ((!sk[1]) & (!g202) & (g358) & (!g360) & (g362) & (!g366)) + ((!sk[1]) & (g202) & (g358) & (!g360) & (g362) & (g366)));
	assign g368 = (((!g11) & (!sk[2]) & (g41) & (!g28) & (!g70)) + ((!g11) & (!sk[2]) & (g41) & (!g28) & (!g70)) + ((!g11) & (!sk[2]) & (!g41) & (g28) & (!g70)) + ((!g11) & (!sk[2]) & (!g41) & (g28) & (g70)));
	assign g369 = (((g50) & (!i_6_) & (!sk[3]) & (!g14) & (!g25) & (!g129)) + ((!g50) & (!i_6_) & (!sk[3]) & (g14) & (!g25) & (!g129)) + ((!g50) & (i_6_) & (!sk[3]) & (!g14) & (g25) & (!g129)) + ((!g50) & (i_6_) & (!sk[3]) & (g14) & (!g25) & (g129)) + ((g50) & (i_6_) & (!sk[3]) & (g14) & (!g25) & (!g129)));
	assign g370 = (((i_6_) & (!g45) & (!sk[4]) & (!g1) & (!g47) & (!g110)) + ((!i_6_) & (!g45) & (!sk[4]) & (g1) & (!g47) & (!g110)) + ((!i_6_) & (g45) & (!sk[4]) & (!g1) & (g47) & (!g110)) + ((i_6_) & (!g45) & (!sk[4]) & (!g1) & (g47) & (g110)) + ((!i_6_) & (!g45) & (sk[4]) & (!g1) & (g47) & (!g110)));
	assign g371 = (((g25) & (!g159) & (!sk[5]) & (!g368) & (!g369) & (!g370)) + ((!g25) & (!g159) & (!sk[5]) & (g368) & (!g369) & (!g370)) + ((!g25) & (g159) & (!sk[5]) & (!g368) & (g369) & (!g370)) + ((g25) & (!g159) & (!sk[5]) & (!g368) & (!g369) & (!g370)) + ((!g25) & (!g159) & (sk[5]) & (!g368) & (!g369) & (!g370)));
	assign g372 = (((i_6_) & (!i_7_) & (!i_8_) & (!g77) & (!sk[6]) & (!g99)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g77) & (!sk[6]) & (!g99)) + ((!i_6_) & (i_7_) & (!i_8_) & (g77) & (!sk[6]) & (!g99)) + ((i_6_) & (!i_7_) & (i_8_) & (g77) & (!sk[6]) & (!g99)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g77) & (!sk[6]) & (g99)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g77) & (sk[6]) & (!g99)));
	assign g373 = (((!g67) & (!g116) & (!sk[7]) & (g290)) + ((!g67) & (!g116) & (sk[7]) & (!g290)) + ((!g67) & (!g116) & (sk[7]) & (!g290)));
	assign g374 = (((!sk[8]) & (g173) & (!g294) & (!g145) & (!g140) & (!g373)) + ((!sk[8]) & (!g173) & (!g294) & (g145) & (!g140) & (!g373)) + ((!sk[8]) & (!g173) & (g294) & (!g145) & (g140) & (!g373)) + ((sk[8]) & (!g173) & (!g294) & (!g145) & (g140) & (g373)));
	assign g375 = (((g23) & (!g75) & (!g160) & (!g372) & (!sk[9]) & (!g374)) + ((!g23) & (!g75) & (g160) & (!g372) & (!sk[9]) & (!g374)) + ((!g23) & (g75) & (!g160) & (g372) & (!sk[9]) & (!g374)) + ((g23) & (!g75) & (!g160) & (!g372) & (!sk[9]) & (g374)) + ((!g23) & (!g75) & (!g160) & (!g372) & (sk[9]) & (g374)));
	assign g376 = (((!sk[10]) & (g50) & (!g35) & (!g1) & (!g12) & (!g184)) + ((!sk[10]) & (!g50) & (!g35) & (g1) & (!g12) & (!g184)) + ((!sk[10]) & (!g50) & (g35) & (!g1) & (g12) & (!g184)) + ((!sk[10]) & (g50) & (!g35) & (!g1) & (g12) & (!g184)) + ((sk[10]) & (!g50) & (g35) & (!g1) & (!g12) & (g184)));
	assign g377 = (((!i_6_) & (!i_7_) & (!i_8_) & (!g24) & (!g64) & (g26)) + ((!i_6_) & (i_7_) & (i_8_) & (!g24) & (g64) & (!g26)));
	assign g378 = (((g204) & (!sk[12]) & (!g376) & (!g246) & (!g249) & (!g377)) + ((!g204) & (!sk[12]) & (!g376) & (g246) & (!g249) & (!g377)) + ((!g204) & (!sk[12]) & (g376) & (!g246) & (g249) & (!g377)) + ((!g204) & (!sk[12]) & (!g376) & (g246) & (g249) & (!g377)));
	assign g379 = (((i_0_) & (!i_1_) & (!sk[13]) & (!i_2_) & (!g23) & (!g123)) + ((!i_0_) & (!i_1_) & (!sk[13]) & (i_2_) & (!g23) & (!g123)) + ((!i_0_) & (i_1_) & (!sk[13]) & (!i_2_) & (g23) & (!g123)) + ((!i_0_) & (!i_1_) & (!sk[13]) & (i_2_) & (!g23) & (g123)) + ((i_0_) & (!i_1_) & (!sk[13]) & (i_2_) & (!g23) & (!g123)));
	assign g380 = (((i_3_) & (!g195) & (!sk[14]) & (!g379) & (!g90) & (!g618)) + ((!i_3_) & (!g195) & (!sk[14]) & (g379) & (!g90) & (!g618)) + ((!i_3_) & (g195) & (!sk[14]) & (!g379) & (g90) & (!g618)) + ((i_3_) & (!g195) & (!sk[14]) & (!g379) & (g90) & (g618)) + ((!i_3_) & (!g195) & (sk[14]) & (!g379) & (g90) & (g618)));
	assign g381 = (((g228) & (g330) & (g371) & (g375) & (g378) & (g380)));
	assign g382 = (((!i_6_) & (g63) & (!g21) & (!g25) & (!g110) & (g218)) + ((!i_6_) & (g63) & (!g21) & (!g25) & (!g110) & (!g218)) + ((i_6_) & (g63) & (!g21) & (!g25) & (g110) & (!g218)));
	assign g383 = (((g27) & (!g45) & (!g6) & (g251) & (g287) & (!g382)) + ((!g27) & (g45) & (!g6) & (g251) & (g287) & (!g382)) + ((!g27) & (!g45) & (!g6) & (g251) & (g287) & (!g382)));
	assign g384 = (((!g27) & (!g42) & (g12) & (!g48) & (!g59) & (!g38)) + ((!g27) & (g42) & (!g12) & (g48) & (!g59) & (!g38)));
	assign g385 = (((g27) & (!g21) & (!g6) & (!sk[19]) & (!g3) & (!g121)) + ((!g27) & (!g21) & (g6) & (!sk[19]) & (!g3) & (!g121)) + ((!g27) & (!g21) & (g6) & (!sk[19]) & (g3) & (!g121)) + ((!g27) & (g21) & (!g6) & (!sk[19]) & (g3) & (!g121)) + ((!g27) & (!g21) & (!g6) & (sk[19]) & (!g3) & (g121)));
	assign g386 = (((!g45) & (g1) & (!g2) & (!g38) & (!g384) & (!g385)) + ((!g45) & (!g1) & (!g2) & (!g38) & (!g384) & (!g385)) + ((g45) & (!g1) & (!g2) & (g38) & (!g384) & (!g385)));
	assign g387 = (((!g63) & (!g42) & (!sk[21]) & (g134)) + ((g63) & (g42) & (!sk[21]) & (g134)));
	assign g388 = (((!sk[22]) & (!g1) & (g159) & (!g150) & (!g387)) + ((!sk[22]) & (!g1) & (!g159) & (g150) & (!g387)) + ((sk[22]) & (!g1) & (!g159) & (!g150) & (!g387)) + ((!sk[22]) & (g1) & (g159) & (!g150) & (!g387)));
	assign g389 = (((!g28) & (g110) & (!sk[23]) & (!g116) & (!g141)) + ((!g28) & (!g110) & (!sk[23]) & (g116) & (!g141)) + ((!g28) & (!g110) & (!sk[23]) & (g116) & (g141)) + ((g28) & (g110) & (!sk[23]) & (g116) & (!g141)));
	assign g390 = (((!g18) & (!sk[24]) & (!g170) & (g389)) + ((!g18) & (sk[24]) & (!g170) & (!g389)));
	assign g391 = (((g127) & (!i_2_) & (!i_6_) & (i_7_) & (!i_8_) & (g3)) + ((g127) & (!i_2_) & (i_6_) & (!i_7_) & (!i_8_) & (g3)));
	assign g392 = (((!i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (!g8) & (!g117)) + ((i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (!g8) & (!g117)) + ((!i_4_) & (i_5_) & (!i_0_) & (i_1_) & (!g8) & (!g117)) + ((!i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (!g8) & (!g117)) + ((!i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (!g8) & (!g117)));
	assign g393 = (((g344) & (!sk[27]) & (!g388) & (!g390) & (!g391) & (!g583)) + ((!g344) & (!sk[27]) & (!g388) & (g390) & (!g391) & (!g583)) + ((!g344) & (!sk[27]) & (g388) & (!g390) & (g391) & (!g583)) + ((!g344) & (!sk[27]) & (g388) & (g390) & (!g391) & (g583)));
	assign g394 = (((g72) & (!g166) & (!sk[28]) & (!g383) & (!g386) & (!g393)) + ((!g72) & (!g166) & (!sk[28]) & (g383) & (!g386) & (!g393)) + ((!g72) & (g166) & (!sk[28]) & (!g383) & (g386) & (!g393)) + ((!g72) & (g166) & (!sk[28]) & (g383) & (g386) & (g393)));
	assign g395 = (((!sk[29]) & (g274) & (!g283) & (!g367) & (!g381) & (!g394)) + ((!sk[29]) & (!g274) & (!g283) & (g367) & (!g381) & (!g394)) + ((!sk[29]) & (!g274) & (g283) & (!g367) & (g381) & (!g394)) + ((!sk[29]) & (g274) & (g283) & (g367) & (g381) & (g394)));
	assign g396 = (((!sk[30]) & (!g8) & (g32) & (!g99) & (!g265)) + ((!sk[30]) & (!g8) & (!g32) & (g99) & (!g265)) + ((!sk[30]) & (g8) & (!g32) & (g99) & (!g265)) + ((!sk[30]) & (!g8) & (g32) & (!g99) & (g265)));
	assign g397 = (((!i_4_) & (g42) & (!sk[31]) & (!g12) & (!g9)) + ((!i_4_) & (!g42) & (!sk[31]) & (g12) & (!g9)) + ((i_4_) & (g42) & (!sk[31]) & (g12) & (!g9)) + ((!i_4_) & (!g42) & (sk[31]) & (!g12) & (g9)));
	assign g398 = (((!sk[32]) & (!i_3_) & (!i_5_) & (g396) & (!g397)) + ((!sk[32]) & (!i_3_) & (i_5_) & (!g396) & (!g397)) + ((sk[32]) & (!i_3_) & (!i_5_) & (!g396) & (!g397)) + ((sk[32]) & (!i_3_) & (!i_5_) & (!g396) & (!g397)));
	assign g399 = (((g21) & (!sk[33]) & (!g42) & (!g12) & (!g75) & (!g124)) + ((!g21) & (!sk[33]) & (!g42) & (g12) & (!g75) & (!g124)) + ((!g21) & (!sk[33]) & (g42) & (!g12) & (g75) & (!g124)) + ((!g21) & (sk[33]) & (!g42) & (!g12) & (!g75) & (!g124)) + ((g21) & (!sk[33]) & (!g42) & (!g12) & (!g75) & (!g124)) + ((!g21) & (!sk[33]) & (!g42) & (g12) & (!g75) & (!g124)));
	assign g400 = (((g2) & (!sk[34]) & (!g3) & (!g9) & (!g243) & (!g399)) + ((!g2) & (!sk[34]) & (!g3) & (g9) & (!g243) & (!g399)) + ((!g2) & (!sk[34]) & (g3) & (!g9) & (g243) & (!g399)) + ((!g2) & (sk[34]) & (!g3) & (!g9) & (!g243) & (g399)) + ((!g2) & (sk[34]) & (!g3) & (!g9) & (!g243) & (g399)) + ((!g2) & (sk[34]) & (!g3) & (!g9) & (!g243) & (g399)) + ((!g2) & (sk[34]) & (!g3) & (!g9) & (!g243) & (g399)));
	assign g401 = (((i_3_) & (!g50) & (!i_0_) & (!i_2_) & (!sk[35]) & (!i_6_)) + ((!i_3_) & (!g50) & (i_0_) & (!i_2_) & (!sk[35]) & (!i_6_)) + ((!i_3_) & (g50) & (!i_0_) & (i_2_) & (!sk[35]) & (!i_6_)) + ((!i_3_) & (g50) & (!i_0_) & (i_2_) & (!sk[35]) & (!i_6_)));
	assign g402 = (((i_6_) & (!sk[36]) & (!g25) & (!g137) & (!g38) & (!g401)) + ((!i_6_) & (!sk[36]) & (!g25) & (g137) & (!g38) & (!g401)) + ((!i_6_) & (!sk[36]) & (!g25) & (g137) & (!g38) & (g401)) + ((!i_6_) & (!sk[36]) & (g25) & (!g137) & (g38) & (!g401)) + ((i_6_) & (!sk[36]) & (!g25) & (g137) & (!g38) & (!g401)));
	assign g403 = (((i_6_) & (i_7_) & (i_8_) & (g77) & (!g71) & (!g161)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g77) & (g71) & (!g161)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g77) & (g71) & (!g161)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g77) & (!g71) & (g161)));
	assign g404 = (((!sk[38]) & (!g402) & (g93) & (!g631) & (!g403)) + ((!sk[38]) & (!g402) & (!g93) & (g631) & (!g403)) + ((!sk[38]) & (!g402) & (g93) & (g631) & (!g403)));
	assign g405 = (((!sk[39]) & (g149) & (!g398) & (!g242) & (!g400) & (!g404)) + ((!sk[39]) & (!g149) & (!g398) & (g242) & (!g400) & (!g404)) + ((!sk[39]) & (!g149) & (g398) & (!g242) & (g400) & (!g404)) + ((!sk[39]) & (!g149) & (g398) & (g242) & (g400) & (g404)));
	assign g406 = (((!i_3_) & (!sk[40]) & (i_0_) & (!i_2_) & (!g85)) + ((!i_3_) & (!sk[40]) & (!i_0_) & (i_2_) & (!g85)) + ((i_3_) & (!sk[40]) & (!i_0_) & (i_2_) & (g85)));
	assign g407 = (((!g50) & (g48) & (g88) & (!sk[41]) & (!g111) & (!g230)) + ((g50) & (!g48) & (!g88) & (!sk[41]) & (!g111) & (!g230)) + ((!g50) & (!g48) & (g88) & (!sk[41]) & (!g111) & (!g230)) + ((!g50) & (g48) & (!g88) & (!sk[41]) & (g111) & (!g230)) + ((g50) & (!g48) & (!g88) & (!sk[41]) & (g111) & (g230)));
	assign g408 = (((g14) & (!g1) & (!g22) & (!sk[42]) & (!g406) & (!g407)) + ((!g14) & (!g1) & (g22) & (!sk[42]) & (!g406) & (!g407)) + ((!g14) & (g1) & (!g22) & (!sk[42]) & (g406) & (!g407)) + ((!g14) & (!g1) & (!g22) & (sk[42]) & (!g406) & (!g407)) + ((!g14) & (g1) & (!g22) & (sk[42]) & (!g406) & (!g407)) + ((!g14) & (g1) & (!g22) & (sk[42]) & (!g406) & (!g407)) + ((!g14) & (!g1) & (!g22) & (sk[42]) & (!g406) & (!g407)));
	assign g409 = (((!i_6_) & (!i_7_) & (i_8_) & (!g33) & (!g184) & (g401)) + ((i_6_) & (i_7_) & (!i_8_) & (g33) & (!g184) & (!g401)) + ((i_6_) & (i_7_) & (i_8_) & (!g33) & (g184) & (!g401)));
	assign g410 = (((!g35) & (g48) & (!g117) & (!sk[44]) & (!g334)) + ((!g35) & (!g48) & (g117) & (!sk[44]) & (!g334)) + ((!g35) & (!g48) & (!g117) & (sk[44]) & (!g334)) + ((!g35) & (!g48) & (!g117) & (sk[44]) & (!g334)));
	assign g411 = (((i_4_) & (!i_5_) & (!i_0_) & (!sk[45]) & (!i_1_) & (!g12)) + ((!i_4_) & (!i_5_) & (i_0_) & (!sk[45]) & (!i_1_) & (!g12)) + ((!i_4_) & (i_5_) & (!i_0_) & (!sk[45]) & (i_1_) & (!g12)) + ((!i_4_) & (!i_5_) & (!i_0_) & (sk[45]) & (i_1_) & (g12)));
	assign g412 = (((g8) & (!g137) & (!g91) & (!sk[46]) & (!g243) & (!g411)) + ((!g8) & (!g137) & (g91) & (!sk[46]) & (!g243) & (!g411)) + ((!g8) & (g137) & (!g91) & (!sk[46]) & (g243) & (!g411)) + ((!g8) & (!g137) & (!g91) & (sk[46]) & (!g243) & (!g411)) + ((!g8) & (!g137) & (!g91) & (sk[46]) & (!g243) & (!g411)) + ((!g8) & (!g137) & (!g91) & (sk[46]) & (!g243) & (!g411)) + ((!g8) & (!g137) & (!g91) & (sk[46]) & (!g243) & (!g411)));
	assign g413 = (((!sk[47]) & (!g2) & (!g70) & (g158)) + ((!sk[47]) & (g2) & (!g70) & (g158)) + ((sk[47]) & (g2) & (g70) & (!g158)));
	assign g414 = (((!sk[48]) & (i_5_) & (!g6) & (!g5) & (!g110) & (!g111)) + ((!sk[48]) & (!i_5_) & (!g6) & (g5) & (!g110) & (!g111)) + ((!sk[48]) & (!i_5_) & (g6) & (!g5) & (g110) & (!g111)) + ((!sk[48]) & (!i_5_) & (g6) & (g5) & (g110) & (!g111)) + ((!sk[48]) & (!i_5_) & (!g6) & (g5) & (g110) & (g111)));
	assign g415 = (((!g23) & (g359) & (!sk[49]) & (!g413) & (!g414)) + ((!g23) & (!g359) & (!sk[49]) & (g413) & (!g414)) + ((!g23) & (!g359) & (sk[49]) & (!g413) & (!g414)) + ((g23) & (!g359) & (sk[49]) & (!g413) & (!g414)));
	assign g416 = (((g87) & (!sk[50]) & (!g346) & (!g410) & (!g412) & (!g415)) + ((!g87) & (!sk[50]) & (!g346) & (g410) & (!g412) & (!g415)) + ((!g87) & (!sk[50]) & (g346) & (!g410) & (g412) & (!g415)) + ((!g87) & (!sk[50]) & (!g346) & (g410) & (g412) & (g415)));
	assign g417 = (((g254) & (!g307) & (!sk[51]) & (!g289) & (!g409) & (!g416)) + ((!g254) & (!g307) & (!sk[51]) & (g289) & (!g409) & (!g416)) + ((!g254) & (g307) & (!sk[51]) & (!g289) & (g409) & (!g416)) + ((g254) & (g307) & (!sk[51]) & (g289) & (!g409) & (g416)));
	assign g418 = (((!g381) & (!sk[52]) & (g405) & (!g408) & (!g417)) + ((!g381) & (!sk[52]) & (!g405) & (g408) & (!g417)) + ((g381) & (!sk[52]) & (g405) & (g408) & (g417)));
	assign g419 = (((i_6_) & (!sk[53]) & (!i_7_) & (!i_8_) & (!g189) & (!g406)) + ((!i_6_) & (!sk[53]) & (!i_7_) & (i_8_) & (!g189) & (!g406)) + ((!i_6_) & (!sk[53]) & (i_7_) & (!i_8_) & (g189) & (!g406)) + ((!i_6_) & (!sk[53]) & (!i_7_) & (i_8_) & (g189) & (!g406)) + ((!i_6_) & (sk[53]) & (i_7_) & (!i_8_) & (!g189) & (g406)));
	assign g420 = (((!i_0_) & (i_1_) & (!i_2_) & (!i_6_) & (!i_7_) & (!i_8_)) + ((!i_0_) & (!i_1_) & (i_2_) & (!i_6_) & (i_7_) & (i_8_)));
	assign g421 = (((!i_0_) & (i_6_) & (!sk[55]) & (!g38) & (!g420)) + ((!i_0_) & (!i_6_) & (!sk[55]) & (g38) & (!g420)) + ((!i_0_) & (!i_6_) & (sk[55]) & (!g38) & (g420)));
	assign g422 = (((g28) & (!sk[56]) & (!g42) & (!g45) & (!g1) & (!g32)) + ((!g28) & (!sk[56]) & (!g42) & (g45) & (!g1) & (!g32)) + ((g28) & (!sk[56]) & (g42) & (!g45) & (!g1) & (!g32)) + ((!g28) & (!sk[56]) & (g42) & (!g45) & (g1) & (!g32)) + ((g28) & (!sk[56]) & (!g42) & (!g45) & (!g1) & (g32)));
	assign g423 = (((g27) & (!g6) & (!g36) & (!g422) & (!sk[57]) & (!g572)) + ((!g27) & (!g6) & (g36) & (!g422) & (!sk[57]) & (!g572)) + ((!g27) & (g6) & (!g36) & (g422) & (!sk[57]) & (!g572)) + ((g27) & (!g6) & (!g36) & (!g422) & (!sk[57]) & (g572)) + ((!g27) & (!g6) & (g36) & (!g422) & (!sk[57]) & (g572)) + ((!g27) & (!g6) & (!g36) & (!g422) & (sk[57]) & (g572)));
	assign g424 = (((g2) & (!sk[58]) & (!g38) & (!g110) & (!g421) & (!g423)) + ((!g2) & (!sk[58]) & (!g38) & (g110) & (!g421) & (!g423)) + ((!g2) & (!sk[58]) & (g38) & (!g110) & (g421) & (!g423)) + ((!g2) & (sk[58]) & (!g38) & (!g110) & (!g421) & (g423)) + ((!g2) & (sk[58]) & (g38) & (!g110) & (!g421) & (g423)) + ((!g2) & (sk[58]) & (!g38) & (!g110) & (!g421) & (g423)));
	assign g425 = (((!sk[59]) & (!i_6_) & (i_8_) & (!g21) & (!g1)) + ((!sk[59]) & (!i_6_) & (!i_8_) & (g21) & (!g1)) + ((sk[59]) & (!i_6_) & (!i_8_) & (!g21) & (!g1)));
	assign g426 = (((!sk[60]) & (!i_6_) & (g14) & (!g32) & (!g110)) + ((!sk[60]) & (!i_6_) & (!g14) & (g32) & (!g110)) + ((!sk[60]) & (i_6_) & (!g14) & (g32) & (g110)) + ((!sk[60]) & (!i_6_) & (g14) & (g32) & (g110)));
	assign g427 = (((!g24) & (g4) & (!g425) & (!sk[61]) & (!g426)) + ((!g24) & (!g4) & (g425) & (!sk[61]) & (!g426)) + ((!g24) & (!g4) & (!g425) & (sk[61]) & (!g426)) + ((g24) & (!g4) & (!g425) & (sk[61]) & (!g426)));
	assign g428 = (((!i_3_) & (!sk[62]) & (i_0_) & (!i_2_) & (!g123)) + ((!i_3_) & (!sk[62]) & (!i_0_) & (i_2_) & (!g123)) + ((!i_3_) & (!sk[62]) & (i_0_) & (i_2_) & (g123)));
	assign g429 = (((!g11) & (!g29) & (!sk[63]) & (g428)) + ((g11) & (!g29) & (sk[63]) & (!g428)) + ((!g11) & (!g29) & (sk[63]) & (!g428)));
	assign g430 = (((!g63) & (!sk[64]) & (g45) & (!g129) & (!g141)) + ((g63) & (!sk[64]) & (!g45) & (g129) & (!g141)) + ((!g63) & (!sk[64]) & (!g45) & (g129) & (!g141)) + ((!g63) & (sk[64]) & (!g45) & (!g129) & (g141)));
	assign g431 = (((!g35) & (!g1) & (g16) & (!sk[65]) & (!g161)) + ((!g35) & (g1) & (!g16) & (!sk[65]) & (!g161)) + ((g35) & (!g1) & (!g16) & (sk[65]) & (g161)));
	assign g432 = (((!i_7_) & (!g8) & (g25) & (!g32) & (!g97) & (!g217)) + ((!i_7_) & (!g8) & (!g25) & (!g32) & (!g97) & (!g217)) + ((!i_7_) & (!g8) & (!g25) & (!g32) & (!g97) & (!g217)) + ((!i_7_) & (!g8) & (!g25) & (!g32) & (!g97) & (!g217)) + ((!i_7_) & (!g8) & (!g25) & (!g32) & (!g97) & (!g217)));
	assign g433 = (((!i_1_) & (g6) & (g33) & (!sk[67]) & (!g38)) + ((!i_1_) & (g6) & (!g33) & (!sk[67]) & (!g38)) + ((!i_1_) & (!g6) & (g33) & (!sk[67]) & (!g38)) + ((i_1_) & (g6) & (!g33) & (!sk[67]) & (!g38)));
	assign g434 = (((!g35) & (!g189) & (!g229) & (!g431) & (g432) & (!g433)) + ((!g35) & (!g189) & (!g229) & (!g431) & (g432) & (!g433)));
	assign g435 = (((g352) & (!g332) & (!g429) & (!g430) & (!sk[69]) & (!g434)) + ((!g352) & (!g332) & (g429) & (!g430) & (!sk[69]) & (!g434)) + ((!g352) & (g332) & (!g429) & (g430) & (!sk[69]) & (!g434)) + ((!g352) & (g332) & (g429) & (!g430) & (!sk[69]) & (g434)));
	assign g436 = (((g419) & (!g367) & (!g424) & (!g427) & (!sk[70]) & (!g435)) + ((!g419) & (!g367) & (g424) & (!g427) & (!sk[70]) & (!g435)) + ((!g419) & (g367) & (!g424) & (g427) & (!sk[70]) & (!g435)) + ((!g419) & (g367) & (g424) & (g427) & (!sk[70]) & (g435)));
	assign g437 = (((g31) & (!sk[71]) & (!g300) & (!g371) & (!g405) & (!g436)) + ((!g31) & (!sk[71]) & (!g300) & (g371) & (!g405) & (!g436)) + ((!g31) & (!sk[71]) & (g300) & (!g371) & (g405) & (!g436)) + ((g31) & (!sk[71]) & (g300) & (g371) & (g405) & (g436)));
	assign g438 = (((!sk[72]) & (!g48) & (!g33) & (g368)) + ((sk[72]) & (!g48) & (!g33) & (!g368)) + ((sk[72]) & (!g48) & (!g33) & (!g368)));
	assign g439 = (((g21) & (!sk[73]) & (!g1) & (!g2) & (!g24) & (!g36)) + ((!g21) & (!sk[73]) & (!g1) & (g2) & (!g24) & (!g36)) + ((!g21) & (!sk[73]) & (g1) & (!g2) & (g24) & (!g36)) + ((!g21) & (!sk[73]) & (!g1) & (g2) & (!g24) & (!g36)) + ((!g21) & (!sk[73]) & (!g1) & (g2) & (!g24) & (!g36)));
	assign g440 = (((!i_3_) & (!i_1_) & (!sk[74]) & (i_2_)) + ((!i_3_) & (!i_1_) & (!sk[74]) & (i_2_)));
	assign g441 = (((!g137) & (!sk[75]) & (!g15) & (g440)) + ((g137) & (!sk[75]) & (g15) & (g440)));
	assign g442 = (((g6) & (!g5) & (!g110) & (!g99) & (!sk[76]) & (!g441)) + ((!g6) & (!g5) & (g110) & (!g99) & (!sk[76]) & (!g441)) + ((!g6) & (g5) & (!g110) & (g99) & (!sk[76]) & (!g441)) + ((!g6) & (!g5) & (!g110) & (!g99) & (sk[76]) & (!g441)) + ((!g6) & (!g5) & (!g110) & (!g99) & (sk[76]) & (!g441)) + ((!g6) & (!g5) & (!g110) & (!g99) & (sk[76]) & (!g441)));
	assign g443 = (((g35) & (!g161) & (!g376) & (!g439) & (!sk[77]) & (!g442)) + ((!g35) & (!g161) & (g376) & (!g439) & (!sk[77]) & (!g442)) + ((!g35) & (g161) & (!g376) & (g439) & (!sk[77]) & (!g442)) + ((!g35) & (!g161) & (!g376) & (!g439) & (sk[77]) & (g442)) + ((!g35) & (!g161) & (!g376) & (!g439) & (sk[77]) & (g442)));
	assign g444 = (((!i_8_) & (g65) & (!sk[78]) & (!g247) & (!g398)) + ((!i_8_) & (!g65) & (!sk[78]) & (g247) & (!g398)) + ((!i_8_) & (!g65) & (sk[78]) & (!g247) & (g398)) + ((!i_8_) & (!g65) & (sk[78]) & (!g247) & (g398)));
	assign g445 = (((g266) & (!g438) & (!sk[79]) & (!g358) & (!g443) & (!g444)) + ((!g266) & (!g438) & (!sk[79]) & (g358) & (!g443) & (!g444)) + ((!g266) & (g438) & (!sk[79]) & (!g358) & (g443) & (!g444)) + ((!g266) & (g438) & (!sk[79]) & (g358) & (g443) & (g444)));
	assign g446 = (((i_3_) & (!i_1_) & (!i_2_) & (!i_7_) & (!sk[80]) & (!g64)) + ((!i_3_) & (!i_1_) & (i_2_) & (!i_7_) & (!sk[80]) & (!g64)) + ((!i_3_) & (i_1_) & (!i_2_) & (i_7_) & (!sk[80]) & (!g64)) + ((i_3_) & (i_1_) & (!i_2_) & (i_7_) & (!sk[80]) & (g64)));
	assign g447 = (((g14) & (!g24) & (!g64) & (!sk[81]) & (!g194) & (!g446)) + ((!g14) & (!g24) & (g64) & (!sk[81]) & (!g194) & (!g446)) + ((!g14) & (g24) & (!g64) & (!sk[81]) & (g194) & (!g446)) + ((!g14) & (g24) & (!g64) & (sk[81]) & (!g194) & (!g446)) + ((!g14) & (!g24) & (!g64) & (sk[81]) & (!g194) & (!g446)) + ((!g14) & (!g24) & (!g64) & (sk[81]) & (!g194) & (!g446)));
	assign g448 = (((!sk[82]) & (!g25) & (!g2) & (g38) & (!g110)) + ((!sk[82]) & (!g25) & (g2) & (!g38) & (!g110)) + ((sk[82]) & (!g25) & (!g2) & (!g38) & (!g110)) + ((!sk[82]) & (g25) & (g2) & (!g38) & (!g110)));
	assign g449 = (((i_5_) & (!sk[83]) & (!g6) & (!g23) & (!g110) & (!g440)) + ((!i_5_) & (!sk[83]) & (!g6) & (g23) & (!g110) & (!g440)) + ((!i_5_) & (!sk[83]) & (!g6) & (g23) & (!g110) & (!g440)) + ((!i_5_) & (!sk[83]) & (g6) & (!g23) & (g110) & (!g440)) + ((!i_5_) & (sk[83]) & (!g6) & (!g23) & (!g110) & (!g440)) + ((!i_5_) & (sk[83]) & (!g6) & (!g23) & (!g110) & (!g440)));
	assign g450 = (((!g255) & (g384) & (!sk[84]) & (!g310) & (!g559)) + ((!g255) & (!g384) & (!sk[84]) & (g310) & (!g559)) + ((!g255) & (!g384) & (!sk[84]) & (g310) & (g559)));
	assign g451 = (((!g50) & (i_6_) & (i_8_) & (g5) & (!g13) & (!g17)) + ((g50) & (!i_6_) & (i_8_) & (!g5) & (!g13) & (g17)));
	assign g452 = (((g275) & (!g402) & (!g670) & (!sk[86]) & (!g147) & (!g451)) + ((!g275) & (!g402) & (g670) & (!sk[86]) & (!g147) & (!g451)) + ((!g275) & (g402) & (!g670) & (!sk[86]) & (g147) & (!g451)) + ((!g275) & (!g402) & (g670) & (!sk[86]) & (g147) & (!g451)));
	assign g453 = (((g80) & (g291) & (g383) & (g427) & (g450) & (g452)));
	assign g454 = (((!sk[88]) & (g109) & (!g341) & (!g408) & (!g445) & (!g453)) + ((!sk[88]) & (!g109) & (!g341) & (g408) & (!g445) & (!g453)) + ((!sk[88]) & (!g109) & (g341) & (!g408) & (g445) & (!g453)) + ((!sk[88]) & (g109) & (g341) & (g408) & (g445) & (g453)));
	assign g455 = (((g127) & (!i_2_) & (!g2) & (!g60) & (!sk[89]) & (!g38)) + ((!g127) & (!i_2_) & (g2) & (!g60) & (!sk[89]) & (!g38)) + ((!g127) & (i_2_) & (!g2) & (g60) & (!sk[89]) & (!g38)) + ((g127) & (!i_2_) & (g2) & (!g60) & (!sk[89]) & (!g38)) + ((g127) & (i_2_) & (!g2) & (g60) & (!sk[89]) & (!g38)));
	assign g456 = (((g23) & (!g66) & (!g189) & (!g455) & (!sk[90]) & (!g315)) + ((!g23) & (!g66) & (g189) & (!g455) & (!sk[90]) & (!g315)) + ((!g23) & (g66) & (!g189) & (g455) & (!sk[90]) & (!g315)) + ((g23) & (!g66) & (!g189) & (!g455) & (!sk[90]) & (!g315)) + ((!g23) & (!g66) & (!g189) & (!g455) & (sk[90]) & (!g315)));
	assign g457 = (((g2) & (!g36) & (!g38) & (!sk[91]) & (!g110) & (!g121)) + ((!g2) & (!g36) & (g38) & (!sk[91]) & (!g110) & (!g121)) + ((g2) & (!g36) & (!g38) & (!sk[91]) & (g110) & (!g121)) + ((!g2) & (g36) & (!g38) & (!sk[91]) & (g110) & (!g121)) + ((!g2) & (!g36) & (!g38) & (sk[91]) & (!g110) & (g121)));
	assign g458 = (((!g63) & (!g64) & (!sk[92]) & (g17)) + ((g63) & (g64) & (!sk[92]) & (g17)));
	assign g459 = (((!g267) & (!g313) & (!g389) & (!g419) & (!g457) & (!g458)));
	assign g460 = (((!i_4_) & (i_5_) & (i_1_) & (i_2_) & (!i_6_) & (g14)) + ((i_4_) & (i_5_) & (!i_1_) & (i_2_) & (i_6_) & (g14)));
	assign g461 = (((!i_3_) & (i_6_) & (!i_8_) & (!sk[95]) & (!g13)) + ((!i_3_) & (!i_6_) & (i_8_) & (!sk[95]) & (!g13)) + ((!i_3_) & (!i_6_) & (!i_8_) & (sk[95]) & (!g13)));
	assign g462 = (((!g27) & (g28) & (!g36) & (!sk[96]) & (!g461)) + ((!g27) & (!g28) & (g36) & (!sk[96]) & (!g461)) + ((!g27) & (!g28) & (g36) & (!sk[96]) & (!g461)) + ((!g27) & (!g28) & (!g36) & (sk[96]) & (!g461)) + ((g27) & (!g28) & (!g36) & (sk[96]) & (!g461)));
	assign g463 = (((i_6_) & (!i_7_) & (!sk[97]) & (!i_8_) & (!g71) & (!g26)) + ((!i_6_) & (!i_7_) & (!sk[97]) & (i_8_) & (!g71) & (!g26)) + ((!i_6_) & (i_7_) & (!sk[97]) & (!i_8_) & (g71) & (!g26)) + ((!i_6_) & (!i_7_) & (!sk[97]) & (i_8_) & (g71) & (!g26)) + ((!i_6_) & (!i_7_) & (sk[97]) & (!i_8_) & (!g71) & (g26)) + ((!i_6_) & (i_7_) & (sk[97]) & (!i_8_) & (!g71) & (g26)));
	assign g464 = (((!g50) & (g47) & (!g94) & (!sk[98]) & (!g401)) + ((!g50) & (!g47) & (g94) & (!sk[98]) & (!g401)) + ((!g50) & (g47) & (!g94) & (!sk[98]) & (g401)) + ((g50) & (g47) & (g94) & (!sk[98]) & (!g401)));
	assign g465 = (((g292) & (!g327) & (!g363) & (!g463) & (!sk[99]) & (!g464)) + ((!g292) & (!g327) & (g363) & (!g463) & (!sk[99]) & (!g464)) + ((!g292) & (g327) & (!g363) & (g463) & (!sk[99]) & (!g464)) + ((!g292) & (g327) & (!g363) & (!g463) & (sk[99]) & (!g464)));
	assign g466 = (((g34) & (!sk[100]) & (!g323) & (!g460) & (!g462) & (!g465)) + ((!g34) & (!sk[100]) & (!g323) & (g460) & (!g462) & (!g465)) + ((!g34) & (!sk[100]) & (g323) & (!g460) & (g462) & (!g465)) + ((!g34) & (!sk[100]) & (g323) & (!g460) & (g462) & (g465)));
	assign g467 = (((g154) & (g216) & (g445) & (g456) & (g459) & (g466)));
	assign g468 = (((!sk[102]) & (!g8) & (g45) & (!g13) & (!g165)) + ((!sk[102]) & (!g8) & (!g45) & (g13) & (!g165)) + ((!sk[102]) & (!g8) & (g45) & (!g13) & (!g165)) + ((!sk[102]) & (!g8) & (!g45) & (g13) & (!g165)) + ((sk[102]) & (!g8) & (!g45) & (!g13) & (!g165)));
	assign g469 = (((g21) & (!g6) & (!g23) & (!sk[103]) & (!g24) & (!g3)) + ((!g21) & (!g6) & (g23) & (!sk[103]) & (!g24) & (!g3)) + ((!g21) & (g6) & (!g23) & (!sk[103]) & (g24) & (!g3)) + ((!g21) & (!g6) & (!g23) & (sk[103]) & (!g24) & (!g3)) + ((!g21) & (g6) & (!g23) & (sk[103]) & (!g24) & (g3)));
	assign g470 = (((g8) & (!g2) & (!sk[104]) & (!g26) & (!g239) & (!g469)) + ((!g8) & (!g2) & (!sk[104]) & (g26) & (!g239) & (!g469)) + ((!g8) & (g2) & (!sk[104]) & (!g26) & (g239) & (!g469)) + ((!g8) & (!g2) & (sk[104]) & (!g26) & (!g239) & (!g469)) + ((!g8) & (!g2) & (!sk[104]) & (g26) & (!g239) & (!g469)));
	assign g471 = (((g102) & (!sk[105]) & (!g208) & (!g278) & (!g40) & (!g470)) + ((!g102) & (!sk[105]) & (!g208) & (g278) & (!g40) & (!g470)) + ((!g102) & (!sk[105]) & (g208) & (!g278) & (g40) & (!g470)) + ((!g102) & (sk[105]) & (!g208) & (!g278) & (g40) & (g470)));
	assign g472 = (((!i_3_) & (!i_0_) & (!sk[106]) & (i_1_)) + ((!i_3_) & (!i_0_) & (sk[106]) & (!i_1_)));
	assign g473 = (((i_4_) & (!i_6_) & (!g4) & (!sk[107]) & (!g110) & (!g472)) + ((!i_4_) & (!i_6_) & (g4) & (!sk[107]) & (!g110) & (!g472)) + ((!i_4_) & (!i_6_) & (g4) & (!sk[107]) & (g110) & (!g472)) + ((!i_4_) & (i_6_) & (!g4) & (!sk[107]) & (g110) & (!g472)) + ((!i_4_) & (!i_6_) & (!g4) & (sk[107]) & (!g110) & (g472)));
	assign g474 = (((!g42) & (g38) & (!sk[108]) & (!g29) & (!g159)) + ((!g42) & (!g38) & (!sk[108]) & (g29) & (!g159)) + ((g42) & (!g38) & (sk[108]) & (!g29) & (g159)));
	assign g475 = (((g694) & (!g473) & (!g400) & (!g409) & (!sk[109]) & (!g474)) + ((!g694) & (!g473) & (g400) & (!g409) & (!sk[109]) & (!g474)) + ((!g694) & (g473) & (!g400) & (g409) & (!sk[109]) & (!g474)) + ((g694) & (!g473) & (g400) & (!g409) & (!sk[109]) & (!g474)));
	assign g476 = (((!sk[110]) & (g36) & (!g121) & (!g468) & (!g471) & (!g475)) + ((!sk[110]) & (!g36) & (!g121) & (g468) & (!g471) & (!g475)) + ((!sk[110]) & (!g36) & (g121) & (!g468) & (g471) & (!g475)) + ((!sk[110]) & (g36) & (!g121) & (g468) & (g471) & (g475)) + ((!sk[110]) & (!g36) & (!g121) & (g468) & (g471) & (g475)));
	assign g477 = (((!g50) & (i_6_) & (!g63) & (!sk[111]) & (!g440)) + ((!g50) & (!i_6_) & (g63) & (!sk[111]) & (!g440)) + ((g50) & (i_6_) & (g63) & (!sk[111]) & (g440)));
	assign g478 = (((!i_6_) & (i_7_) & (i_8_) & (g181) & (!g105) & (!g359)) + ((i_6_) & (!i_7_) & (!i_8_) & (g181) & (!g105) & (!g359)) + ((i_6_) & (!i_7_) & (i_8_) & (!g181) & (!g105) & (!g359)) + ((i_6_) & (i_7_) & (!i_8_) & (!g181) & (!g105) & (g359)));
	assign g479 = (((g41) & (!sk[113]) & (!g32) & (!g343) & (!g549) & (!g478)) + ((!g41) & (!sk[113]) & (!g32) & (g343) & (!g549) & (!g478)) + ((!g41) & (!sk[113]) & (g32) & (!g343) & (g549) & (!g478)) + ((!g41) & (!sk[113]) & (!g32) & (g343) & (g549) & (!g478)) + ((!g41) & (!sk[113]) & (!g32) & (g343) & (g549) & (!g478)));
	assign g480 = (((g43) & (!sk[114]) & (!g92) & (!g257) & (!g477) & (!g479)) + ((!g43) & (!sk[114]) & (!g92) & (g257) & (!g477) & (!g479)) + ((!g43) & (!sk[114]) & (g92) & (!g257) & (g477) & (!g479)) + ((!g43) & (!sk[114]) & (!g92) & (g257) & (!g477) & (g479)));
	assign g481 = (((g46) & (!g60) & (!g226) & (!g396) & (!sk[115]) & (!g456)) + ((!g46) & (!g60) & (g226) & (!g396) & (!sk[115]) & (!g456)) + ((!g46) & (g60) & (!g226) & (g396) & (!sk[115]) & (!g456)) + ((!g46) & (!g60) & (!g226) & (!g396) & (sk[115]) & (g456)) + ((!g46) & (!g60) & (!g226) & (!g396) & (sk[115]) & (g456)));
	assign g482 = (((g101) & (!sk[116]) & (!g152) & (!g424) & (!g480) & (!g481)) + ((!g101) & (!sk[116]) & (!g152) & (g424) & (!g480) & (!g481)) + ((!g101) & (!sk[116]) & (g152) & (!g424) & (g480) & (!g481)) + ((!g101) & (!sk[116]) & (g152) & (g424) & (g480) & (g481)));
	assign g483 = (((g21) & (!g12) & (!sk[117]) & (!g6) & (!g13) & (!g110)) + ((!g21) & (!g12) & (!sk[117]) & (g6) & (!g13) & (!g110)) + ((!g21) & (g12) & (!sk[117]) & (!g6) & (g13) & (!g110)) + ((!g21) & (!g12) & (!sk[117]) & (g6) & (!g13) & (g110)) + ((!g21) & (g12) & (sk[117]) & (!g6) & (!g13) & (!g110)));
	assign g484 = (((g28) & (!g25) & (!g12) & (!g32) & (!sk[118]) & (!g36)) + ((!g28) & (!g25) & (g12) & (!g32) & (!sk[118]) & (!g36)) + ((!g28) & (!g25) & (g12) & (g32) & (!sk[118]) & (!g36)) + ((!g28) & (g25) & (!g12) & (g32) & (!sk[118]) & (!g36)) + ((g28) & (!g25) & (!g12) & (!g32) & (!sk[118]) & (!g36)));
	assign g485 = (((!g11) & (!g27) & (!g45) & (!g48) & (g2) & (!g24)) + ((!g11) & (!g27) & (!g45) & (g48) & (!g2) & (!g24)) + ((!g11) & (!g27) & (!g45) & (!g48) & (g2) & (!g24)));
	assign g486 = (((!g1) & (g6) & (!g23) & (!g3) & (g49) & (!g110)) + ((!g1) & (!g6) & (!g23) & (g3) & (!g49) & (!g110)) + ((!g1) & (g6) & (!g23) & (g3) & (!g49) & (g110)));
	assign g487 = (((g155) & (!g483) & (!g484) & (!g485) & (!sk[121]) & (!g486)) + ((!g155) & (!g483) & (g484) & (!g485) & (!sk[121]) & (!g486)) + ((!g155) & (g483) & (!g484) & (g485) & (!sk[121]) & (!g486)) + ((!g155) & (!g483) & (!g484) & (!g485) & (sk[121]) & (!g486)));
	assign g488 = (((!i_6_) & (i_7_) & (!g188) & (!sk[122]) & (!g129)) + ((!i_6_) & (!i_7_) & (g188) & (!sk[122]) & (!g129)) + ((!i_6_) & (!i_7_) & (!g188) & (sk[122]) & (!g129)) + ((!i_6_) & (!i_7_) & (!g188) & (sk[122]) & (!g129)));
	assign g489 = (((i_6_) & (!g32) & (!g18) & (!sk[123]) & (!g110) & (!g488)) + ((!i_6_) & (!g32) & (g18) & (!sk[123]) & (!g110) & (!g488)) + ((!i_6_) & (g32) & (!g18) & (!sk[123]) & (g110) & (!g488)) + ((!i_6_) & (!g32) & (!g18) & (sk[123]) & (!g110) & (g488)) + ((!i_6_) & (!g32) & (!g18) & (sk[123]) & (!g110) & (g488)) + ((!i_6_) & (!g32) & (!g18) & (sk[123]) & (!g110) & (g488)));
	assign g490 = (((!g476) & (g482) & (!g487) & (!sk[124]) & (!g489)) + ((!g476) & (!g482) & (g487) & (!sk[124]) & (!g489)) + ((g476) & (g482) & (g487) & (!sk[124]) & (g489)));
	assign g491 = (((!i_5_) & (!g48) & (!sk[125]) & (g472)) + ((!i_5_) & (g48) & (!sk[125]) & (g472)));
	assign g492 = (((!g1) & (!sk[126]) & (g12) & (!g3) & (!g290)) + ((!g1) & (!sk[126]) & (!g12) & (g3) & (!g290)) + ((g1) & (sk[126]) & (!g12) & (!g3) & (!g290)) + ((!g1) & (sk[126]) & (!g12) & (!g3) & (!g290)) + ((!g1) & (sk[126]) & (!g12) & (!g3) & (!g290)));
	assign g493 = (((g11) & (!g41) & (g45) & (!g29) & (!sk[127]) & (!g141)) + ((g11) & (!g41) & (!g45) & (!g29) & (!sk[127]) & (!g141)) + ((!g11) & (!g41) & (g45) & (!g29) & (!sk[127]) & (!g141)) + ((!g11) & (!g41) & (g45) & (!g29) & (!sk[127]) & (!g141)) + ((g11) & (!g41) & (!g45) & (!g29) & (!sk[127]) & (!g141)) + ((!g11) & (g41) & (!g45) & (g29) & (!sk[127]) & (!g141)) + ((!g11) & (!g41) & (!g45) & (!g29) & (sk[127]) & (!g141)));
	assign g494 = (((g21) & (!g48) & (!g49) & (!sk[0]) & (!g110) & (!g364)) + ((!g21) & (!g48) & (g49) & (!sk[0]) & (!g110) & (!g364)) + ((!g21) & (g48) & (!g49) & (!sk[0]) & (g110) & (!g364)) + ((g21) & (!g48) & (!g49) & (!sk[0]) & (!g110) & (!g364)) + ((!g21) & (!g48) & (!g49) & (sk[0]) & (!g110) & (!g364)) + ((!g21) & (!g48) & (!g49) & (sk[0]) & (!g110) & (!g364)));
	assign g495 = (((g23) & (!g184) & (!sk[1]) & (!g492) & (!g493) & (!g494)) + ((!g23) & (!g184) & (!sk[1]) & (g492) & (!g493) & (!g494)) + ((!g23) & (g184) & (!sk[1]) & (!g492) & (g493) & (!g494)) + ((g23) & (!g184) & (!sk[1]) & (g492) & (g493) & (g494)) + ((!g23) & (!g184) & (!sk[1]) & (g492) & (g493) & (g494)));
	assign g496 = (((g23) & (!g91) & (!g296) & (!g491) & (!sk[2]) & (!g495)) + ((!g23) & (!g91) & (g296) & (!g491) & (!sk[2]) & (!g495)) + ((!g23) & (g91) & (!g296) & (g491) & (!sk[2]) & (!g495)) + ((g23) & (!g91) & (!g296) & (!g491) & (!sk[2]) & (g495)) + ((!g23) & (!g91) & (!g296) & (!g491) & (sk[2]) & (g495)));
	assign g497 = (((g11) & (!sk[3]) & (!i_6_) & (!g2) & (!g32) & (!g110)) + ((!g11) & (!sk[3]) & (!i_6_) & (g2) & (!g32) & (!g110)) + ((!g11) & (!sk[3]) & (i_6_) & (!g2) & (g32) & (!g110)) + ((!g11) & (!sk[3]) & (!i_6_) & (g2) & (!g32) & (g110)) + ((!g11) & (!sk[3]) & (i_6_) & (!g2) & (g32) & (g110)));
	assign g498 = (((!sk[4]) & (g35) & (!g74) & (!g189) & (!g359) & (!g497)) + ((!sk[4]) & (!g35) & (!g74) & (g189) & (!g359) & (!g497)) + ((!sk[4]) & (!g35) & (g74) & (!g189) & (g359) & (!g497)) + ((sk[4]) & (!g35) & (!g74) & (!g189) & (!g359) & (!g497)) + ((!sk[4]) & (g35) & (!g74) & (!g189) & (!g359) & (!g497)));
	assign g499 = (((!i_0_) & (i_1_) & (!i_2_) & (!sk[5]) & (!g194)) + ((!i_0_) & (!i_1_) & (i_2_) & (!sk[5]) & (!g194)) + ((!i_0_) & (!i_1_) & (!i_2_) & (sk[5]) & (!g194)) + ((!i_0_) & (!i_1_) & (!i_2_) & (sk[5]) & (g194)));
	assign g500 = (((g35) & (!g25) & (!sk[6]) & (!g22) & (!g36) & (!g499)) + ((!g35) & (!g25) & (!sk[6]) & (g22) & (!g36) & (!g499)) + ((!g35) & (g25) & (!sk[6]) & (!g22) & (g36) & (!g499)) + ((!g35) & (!g25) & (sk[6]) & (!g22) & (!g36) & (!g499)) + ((!g35) & (g25) & (sk[6]) & (!g22) & (!g36) & (!g499)) + ((!g35) & (!g25) & (sk[6]) & (!g22) & (g36) & (!g499)));
	assign g501 = (((g23) & (!g71) & (!g294) & (!sk[7]) & (!g88) & (!g212)) + ((!g23) & (!g71) & (g294) & (!sk[7]) & (!g88) & (!g212)) + ((!g23) & (g71) & (!g294) & (!sk[7]) & (g88) & (!g212)) + ((g23) & (!g71) & (!g294) & (!sk[7]) & (!g88) & (!g212)) + ((!g23) & (!g71) & (!g294) & (sk[7]) & (!g88) & (!g212)));
	assign g502 = (((g27) & (!g12) & (!sk[8]) & (!g33) & (!g4) & (!g194)) + ((!g27) & (!g12) & (!sk[8]) & (g33) & (!g4) & (!g194)) + ((g27) & (!g12) & (!sk[8]) & (!g33) & (!g4) & (!g194)) + ((!g27) & (g12) & (!sk[8]) & (!g33) & (g4) & (!g194)) + ((!g27) & (!g12) & (sk[8]) & (!g33) & (!g4) & (!g194)) + ((!g27) & (!g12) & (!sk[8]) & (g33) & (!g4) & (!g194)));
	assign g503 = (((!sk[9]) & (g174) & (!g277) & (!g500) & (!g501) & (!g502)) + ((!sk[9]) & (!g174) & (!g277) & (g500) & (!g501) & (!g502)) + ((!sk[9]) & (!g174) & (g277) & (!g500) & (g501) & (!g502)) + ((!sk[9]) & (!g174) & (!g277) & (g500) & (g501) & (g502)));
	assign g504 = (((!g6) & (!sk[10]) & (g59) & (!g88) & (!g265)) + ((g6) & (!sk[10]) & (!g59) & (g88) & (!g265)) + ((!g6) & (!sk[10]) & (!g59) & (g88) & (!g265)) + ((!g6) & (sk[10]) & (!g59) & (!g88) & (g265)));
	assign g505 = (((!g37) & (g129) & (!g386) & (!sk[11]) & (!g504)) + ((!g37) & (!g129) & (g386) & (!sk[11]) & (!g504)) + ((!g37) & (!g129) & (g386) & (!sk[11]) & (!g504)) + ((!g37) & (!g129) & (g386) & (!sk[11]) & (!g504)));
	assign g506 = (((!sk[12]) & (g179) & (!g438) & (!g498) & (!g503) & (!g505)) + ((!sk[12]) & (!g179) & (!g438) & (g498) & (!g503) & (!g505)) + ((!sk[12]) & (!g179) & (g438) & (!g498) & (g503) & (!g505)) + ((!sk[12]) & (!g179) & (g438) & (g498) & (g503) & (g505)));
	assign g507 = (((!sk[13]) & (!g35) & (!g45) & (g13)) + ((sk[13]) & (g35) & (!g45) & (!g13)));
	assign g508 = (((i_3_) & (!sk[14]) & (!g50) & (!g127) & (!g8) & (!g84)) + ((!i_3_) & (!sk[14]) & (!g50) & (g127) & (!g8) & (!g84)) + ((!i_3_) & (!sk[14]) & (g50) & (!g127) & (g8) & (!g84)) + ((!i_3_) & (sk[14]) & (!g50) & (!g127) & (g8) & (g84)) + ((!i_3_) & (!sk[14]) & (g50) & (g127) & (g8) & (!g84)));
	assign g509 = (((g63) & (!sk[15]) & (!g6) & (!g129) & (!g507) & (!g508)) + ((!g63) & (!sk[15]) & (!g6) & (g129) & (!g507) & (!g508)) + ((!g63) & (!sk[15]) & (g6) & (!g129) & (g507) & (!g508)) + ((!g63) & (sk[15]) & (!g6) & (!g129) & (!g507) & (!g508)) + ((!g63) & (!sk[15]) & (!g6) & (g129) & (!g507) & (!g508)));
	assign g510 = (((!g476) & (g496) & (!g506) & (!sk[16]) & (!g509)) + ((!g476) & (!g496) & (g506) & (!sk[16]) & (!g509)) + ((g476) & (g496) & (g506) & (!sk[16]) & (g509)));
	assign g511 = (((!g21) & (!g25) & (g48) & (!g2) & (!g13) & (!g38)) + ((!g21) & (!g25) & (!g48) & (g2) & (!g13) & (!g38)) + ((!g21) & (!g25) & (!g48) & (g2) & (!g13) & (!g38)));
	assign g512 = (((!g42) & (g12) & (!sk[18]) & (!g59) & (!g7)) + ((!g42) & (!g12) & (!sk[18]) & (g59) & (!g7)) + ((g42) & (g12) & (!sk[18]) & (!g59) & (!g7)) + ((!g42) & (!g12) & (sk[18]) & (!g59) & (g7)));
	assign g513 = (((!g27) & (!sk[19]) & (g45) & (!g23) & (!g512)) + ((!g27) & (!sk[19]) & (!g45) & (g23) & (!g512)) + ((!g27) & (!sk[19]) & (g45) & (!g23) & (!g512)) + ((!g27) & (!sk[19]) & (!g45) & (g23) & (!g512)) + ((g27) & (sk[19]) & (!g45) & (!g23) & (!g512)));
	assign g514 = (((g41) & (!g21) & (!g3) & (!sk[20]) & (!g29) & (!g265)) + ((!g41) & (!g21) & (g3) & (!sk[20]) & (!g29) & (!g265)) + ((!g41) & (g21) & (!g3) & (sk[20]) & (!g29) & (!g265)) + ((!g41) & (!g21) & (!g3) & (sk[20]) & (!g29) & (!g265)) + ((!g41) & (g21) & (!g3) & (!sk[20]) & (g29) & (!g265)) + ((!g41) & (!g21) & (!g3) & (sk[20]) & (!g29) & (!g265)));
	assign g515 = (((g134) & (!g413) & (!g457) & (!g472) & (!sk[21]) & (!g514)) + ((!g134) & (!g413) & (g457) & (!g472) & (!sk[21]) & (!g514)) + ((!g134) & (g413) & (!g457) & (g472) & (!sk[21]) & (!g514)) + ((!g134) & (!g413) & (!g457) & (!g472) & (sk[21]) & (g514)) + ((!g134) & (!g413) & (!g457) & (!g472) & (sk[21]) & (g514)));
	assign g516 = (((!g28) & (g32) & (g67) & (!sk[22]) & (!g181)) + ((!g28) & (g32) & (!g67) & (!sk[22]) & (!g181)) + ((!g28) & (!g32) & (g67) & (!sk[22]) & (!g181)) + ((g28) & (!g32) & (!g67) & (sk[22]) & (g181)));
	assign g517 = (((!g314) & (g293) & (!sk[23]) & (!g236) & (!g516)) + ((!g314) & (!g293) & (!sk[23]) & (g236) & (!g516)) + ((!g314) & (!g293) & (!sk[23]) & (g236) & (!g516)));
	assign g518 = (((!sk[24]) & (g122) & (!g511) & (!g513) & (!g543) & (!g517)) + ((!sk[24]) & (!g122) & (!g511) & (g513) & (!g543) & (!g517)) + ((!sk[24]) & (!g122) & (g511) & (!g513) & (g543) & (!g517)) + ((!sk[24]) & (!g122) & (!g511) & (g513) & (g543) & (g517)));
	assign g519 = (((!g13) & (!sk[25]) & (g123) & (!g387) & (!g458)) + ((!g13) & (!sk[25]) & (!g123) & (g387) & (!g458)) + ((!g13) & (sk[25]) & (!g123) & (!g387) & (!g458)) + ((g13) & (!sk[25]) & (g123) & (!g387) & (!g458)));
	assign g520 = (((g431) & (!sk[26]) & (!g487) & (!g506) & (!g518) & (!g519)) + ((!g431) & (!sk[26]) & (!g487) & (g506) & (!g518) & (!g519)) + ((!g431) & (!sk[26]) & (g487) & (!g506) & (g518) & (!g519)) + ((!g431) & (!sk[26]) & (g487) & (g506) & (g518) & (g519)));
	assign g521 = (((!sk[27]) & (!g8) & (!g117) & (g428)) + ((sk[27]) & (!g8) & (!g117) & (!g428)) + ((sk[27]) & (!g8) & (!g117) & (!g428)));
	assign g522 = (((!i_4_) & (!i_5_) & (!g63) & (!g65) & (!g472) & (g521)) + ((i_4_) & (!i_5_) & (!g63) & (!g65) & (!g472) & (g521)) + ((!i_4_) & (i_5_) & (!g63) & (!g65) & (!g472) & (g521)) + ((!i_4_) & (!i_5_) & (!g63) & (!g65) & (!g472) & (g521)));
	assign g523 = (((!g482) & (g496) & (!g518) & (!sk[29]) & (!g522)) + ((!g482) & (!g496) & (g518) & (!sk[29]) & (!g522)) + ((g482) & (g496) & (g518) & (!sk[29]) & (g522)));
	assign g524 = (((g28) & (!g25) & (!sk[30]) & (!g38) & (!g110) & (!g159)) + ((!g28) & (!g25) & (!sk[30]) & (g38) & (!g110) & (!g159)) + ((g28) & (!g25) & (!sk[30]) & (!g38) & (!g110) & (!g159)) + ((!g28) & (g25) & (!sk[30]) & (!g38) & (g110) & (!g159)) + ((!g28) & (!g25) & (sk[30]) & (!g38) & (g110) & (g159)));
	assign g525 = (((i_6_) & (!i_7_) & (!i_8_) & (!g45) & (!g3) & (g110)) + ((i_6_) & (i_7_) & (!i_8_) & (!g45) & (g3) & (g110)));
	assign g526 = (((!i_6_) & (i_7_) & (!i_8_) & (!g21) & (!g25) & (!g110)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g21) & (!g25) & (g110)));
	assign g527 = (((i_6_) & (!sk[33]) & (!i_7_) & (!i_8_) & (!g46) & (!g184)) + ((!i_6_) & (!sk[33]) & (!i_7_) & (i_8_) & (!g46) & (!g184)) + ((!i_6_) & (!sk[33]) & (i_7_) & (!i_8_) & (g46) & (!g184)) + ((!i_6_) & (sk[33]) & (!i_7_) & (!i_8_) & (!g46) & (g184)) + ((!i_6_) & (sk[33]) & (!i_7_) & (!i_8_) & (g46) & (!g184)) + ((!i_6_) & (!sk[33]) & (!i_7_) & (i_8_) & (!g46) & (g184)));
	assign g528 = (((!g500) & (g525) & (!g526) & (!sk[34]) & (!g527)) + ((!g500) & (!g525) & (g526) & (!sk[34]) & (!g527)) + ((g500) & (!g525) & (!g526) & (sk[34]) & (!g527)));
	assign g529 = (((i_6_) & (!i_7_) & (!sk[35]) & (!i_8_) & (!g189) & (!g161)) + ((!i_6_) & (!i_7_) & (!sk[35]) & (i_8_) & (!g189) & (!g161)) + ((!i_6_) & (i_7_) & (!sk[35]) & (!i_8_) & (g189) & (!g161)) + ((i_6_) & (i_7_) & (!sk[35]) & (!i_8_) & (!g189) & (g161)) + ((i_6_) & (!i_7_) & (!sk[35]) & (i_8_) & (!g189) & (g161)) + ((i_6_) & (!i_7_) & (!sk[35]) & (i_8_) & (g189) & (!g161)));
	assign g530 = (((!g25) & (g23) & (!g38) & (!sk[36]) & (!g491)) + ((!g25) & (!g23) & (g38) & (!sk[36]) & (!g491)) + ((!g25) & (g23) & (!g38) & (!sk[36]) & (!g491)) + ((!g25) & (!g23) & (g38) & (!sk[36]) & (!g491)) + ((g25) & (!g23) & (!g38) & (sk[36]) & (!g491)));
	assign g531 = (((!g473) & (g498) & (!g529) & (!sk[37]) & (!g530)) + ((!g473) & (!g498) & (g529) & (!sk[37]) & (!g530)) + ((!g473) & (g498) & (!g529) & (!sk[37]) & (g530)));
	assign g532 = (((!g524) & (!g528) & (!sk[38]) & (g531)) + ((!g524) & (g528) & (!sk[38]) & (g531)));
	assign g533 = (((g35) & (!g23) & (!g36) & (!g110) & (!sk[39]) & (!g99)) + ((!g35) & (!g23) & (g36) & (!g110) & (!sk[39]) & (!g99)) + ((g35) & (!g23) & (!g36) & (g110) & (!sk[39]) & (!g99)) + ((!g35) & (g23) & (!g36) & (g110) & (!sk[39]) & (!g99)) + ((!g35) & (!g23) & (!g36) & (!g110) & (sk[39]) & (g99)));
	assign g534 = (((i_0_) & (!i_1_) & (!i_2_) & (!sk[40]) & (!g2) & (!g59)) + ((!i_0_) & (!i_1_) & (i_2_) & (!sk[40]) & (!g2) & (!g59)) + ((!i_0_) & (i_1_) & (!i_2_) & (!sk[40]) & (g2) & (!g59)) + ((!i_0_) & (!i_1_) & (!i_2_) & (sk[40]) & (!g2) & (!g59)) + ((!i_0_) & (!i_1_) & (!i_2_) & (sk[40]) & (g2) & (!g59)));
	assign g535 = (((!g6) & (g23) & (!sk[41]) & (!g189) & (!g99)) + ((!g6) & (!g23) & (!sk[41]) & (g189) & (!g99)) + ((g6) & (!g23) & (sk[41]) & (!g189) & (g99)));
	assign g536 = (((g28) & (!g38) & (!sk[42]) & (!g110) & (!g534) & (!g535)) + ((!g28) & (!g38) & (!sk[42]) & (g110) & (!g534) & (!g535)) + ((!g28) & (g38) & (!sk[42]) & (!g110) & (g534) & (!g535)) + ((!g28) & (!g38) & (sk[42]) & (!g110) & (!g534) & (!g535)) + ((!g28) & (g38) & (sk[42]) & (!g110) & (!g534) & (!g535)) + ((!g28) & (!g38) & (sk[42]) & (!g110) & (!g534) & (!g535)));
	assign g537 = (((!g533) & (!g531) & (!sk[43]) & (g536)) + ((!g533) & (g531) & (!sk[43]) & (g536)));
	assign g538 = (((g8) & (g46) & (!sk[44]) & (!g2) & (!g26)) + ((!g8) & (g46) & (!sk[44]) & (!g2) & (!g26)) + ((!g8) & (!g46) & (!sk[44]) & (g2) & (!g26)) + ((!g8) & (!g46) & (!sk[44]) & (g2) & (g26)));
	assign g539 = (((!sk[45]) & (i_4_) & (!i_6_) & (!g6) & (!g161) & (!g472)) + ((!sk[45]) & (!i_4_) & (!i_6_) & (g6) & (!g161) & (!g472)) + ((!sk[45]) & (!i_4_) & (!i_6_) & (g6) & (g161) & (!g472)) + ((!sk[45]) & (!i_4_) & (i_6_) & (!g6) & (g161) & (!g472)) + ((sk[45]) & (!i_4_) & (!i_6_) & (!g6) & (!g161) & (g472)));
	assign g540 = (((g497) & (!g524) & (!g538) & (!g536) & (!sk[46]) & (!g539)) + ((!g497) & (!g524) & (g538) & (!g536) & (!sk[46]) & (!g539)) + ((!g497) & (g524) & (!g538) & (g536) & (!sk[46]) & (!g539)) + ((!g497) & (!g524) & (!g538) & (g536) & (sk[46]) & (!g539)));
	assign g541 = (((i_4_) & (!sk[47]) & (!i_5_) & (!i_6_) & (!g63) & (!g472)) + ((!i_4_) & (!sk[47]) & (!i_5_) & (i_6_) & (!g63) & (!g472)) + ((!i_4_) & (!sk[47]) & (i_5_) & (!i_6_) & (g63) & (!g472)) + ((!i_4_) & (sk[47]) & (!i_5_) & (!i_6_) & (!g63) & (g472)) + ((!i_4_) & (!sk[47]) & (!i_5_) & (i_6_) & (g63) & (g472)));
	assign g542 = (((!g533) & (g538) & (!sk[48]) & (!g541) & (!g528)) + ((!g533) & (!g538) & (!sk[48]) & (g541) & (!g528)) + ((!g533) & (!g538) & (sk[48]) & (!g541) & (g528)));
	assign g543 = (((g515) & (!sk[49]) & (g544)) + ((!g515) & (!sk[49]) & (g544)));
	assign g544 = (((!sk[50]) & (!g545) & (g546)) + ((sk[50]) & (!g545) & (!g546)));
	assign g545 = (((!i_6_) & (!sk[51]) & (g547)) + ((!i_6_) & (!sk[51]) & (g547)));
	assign g546 = (((i_6_) & (!sk[52]) & (g548)) + ((!i_6_) & (!sk[52]) & (g548)));
	assign g547 = (((!i_8_) & (!g88) & (sk[53]) & (!i_7_)) + ((i_8_) & (!g88) & (!sk[53]) & (i_7_)) + ((!i_8_) & (!g88) & (!sk[53]) & (i_7_)) + ((!i_8_) & (!g88) & (sk[53]) & (!i_7_)));
	assign g548 = (((!g98) & (i_8_) & (!sk[54]) & (!g73) & (!i_7_)) + ((!g98) & (!i_8_) & (!sk[54]) & (g73) & (!i_7_)) + ((!g98) & (!i_8_) & (sk[54]) & (!g73) & (!i_7_)) + ((!g98) & (!i_8_) & (sk[54]) & (!g73) & (!i_7_)));
	assign g549 = (((!sk[55]) & (!g550) & (g551)) + ((sk[55]) & (!g550) & (!g551)));
	assign g550 = (((!sk[56]) & (!i_0_) & (g552)) + ((!sk[56]) & (!i_0_) & (g552)));
	assign g551 = (((i_0_) & (!sk[57]) & (g554)) + ((!i_0_) & (!sk[57]) & (g554)));
	assign g552 = (((!sk[58]) & (!i_1_) & (g553)) + ((sk[58]) & (!i_1_) & (!g553)));
	assign g553 = (((!i_1_) & (!sk[59]) & (i_2_)) + ((!i_1_) & (!sk[59]) & (i_2_)));
	assign g554 = (((!g555) & (!sk[60]) & (g556)) + ((!g555) & (sk[60]) & (!g556)));
	assign g555 = (((!i_1_) & (!sk[61]) & (g557)) + ((!i_1_) & (!sk[61]) & (g557)));
	assign g556 = (((i_1_) & (!sk[62]) & (g558)) + ((!i_1_) & (!sk[62]) & (g558)));
	assign g557 = (((!g36) & (g23) & (!g6) & (!sk[63]) & (!i_2_)) + ((g36) & (!g23) & (!g6) & (sk[63]) & (!i_2_)) + ((!g36) & (!g23) & (g6) & (!sk[63]) & (!i_2_)) + ((!g36) & (!g23) & (!g6) & (sk[63]) & (i_2_)));
	assign g558 = (((!g16) & (!sk[64]) & (i_2_)) + ((!g16) & (sk[64]) & (!i_2_)));
	assign g559 = (((!sk[65]) & (!g560) & (g561)) + ((sk[65]) & (!g560) & (!g561)));
	assign g560 = (((!sk[66]) & (!g243) & (g562)) + ((!sk[66]) & (!g243) & (g562)));
	assign g561 = (((!sk[67]) & (!g243) & (g565)) + ((!sk[67]) & (g243) & (g565)));
	assign g562 = (((!sk[68]) & (!g563) & (g564)) + ((sk[68]) & (!g563) & (!g564)));
	assign g563 = (((!i_8_) & (!sk[69]) & (g568)) + ((!i_8_) & (!sk[69]) & (g568)));
	assign g564 = (((i_8_) & (!sk[70]) & (g569)) + ((!i_8_) & (!sk[70]) & (g569)));
	assign g565 = (((!sk[71]) & (!g566) & (g567)) + ((sk[71]) & (!g566) & (!g567)));
	assign g566 = (((!sk[72]) & (!i_8_) & (g570)) + ((!sk[72]) & (!i_8_) & (g570)));
	assign g567 = (((!sk[73]) & (!i_8_) & (g571)) + ((!sk[73]) & (i_8_) & (g571)));
	assign g568 = (((!g448) & (!sk[74]) & (!g449) & (g447)) + ((g448) & (!sk[74]) & (g449) & (g447)));
	assign g569 = (((!g448) & (!sk[75]) & (!g449) & (g447)) + ((g448) & (!sk[75]) & (g449) & (g447)));
	assign g570 = (((!sk[76]) & (!g448) & (g449) & (!i_7_) & (!g447)) + ((!sk[76]) & (!g448) & (!g449) & (i_7_) & (!g447)) + ((!sk[76]) & (g448) & (g449) & (i_7_) & (g447)));
	assign g571 = (((!g448) & (!sk[77]) & (g449) & (!i_6_) & (!g447)) + ((!g448) & (!sk[77]) & (!g449) & (i_6_) & (!g447)) + ((g448) & (!sk[77]) & (g449) & (i_6_) & (g447)));
	assign g572 = (((!sk[78]) & (!g573) & (g574)) + ((sk[78]) & (!g573) & (!g574)));
	assign g573 = (((!i_6_) & (!sk[79]) & (g575)) + ((!i_6_) & (!sk[79]) & (g575)));
	assign g574 = (((!sk[80]) & (!i_6_) & (g578)) + ((!sk[80]) & (i_6_) & (g578)));
	assign g575 = (((!sk[81]) & (!g576) & (g577)) + ((sk[81]) & (!g576) & (!g577)));
	assign g576 = (((!i_8_) & (!sk[82]) & (g580)) + ((!i_8_) & (!sk[82]) & (g580)));
	assign g577 = (((i_8_) & (!sk[83]) & (g581)) + ((!i_8_) & (!sk[83]) & (g581)));
	assign g578 = (((!i_8_) & (!sk[84]) & (g579)) + ((!i_8_) & (sk[84]) & (!g579)));
	assign g579 = (((!sk[85]) & (!i_8_) & (g582)) + ((!sk[85]) & (!i_8_) & (g582)));
	assign g580 = (((!sk[86]) & (!g59) & (!g25) & (i_7_)) + ((sk[86]) & (g59) & (!g25) & (!i_7_)) + ((sk[86]) & (!g59) & (g25) & (!i_7_)));
	assign g581 = (((!g59) & (!sk[87]) & (g13)) + ((g59) & (sk[87]) & (!g13)));
	assign g582 = (((!i_7_) & (!sk[88]) & (g105)) + ((i_7_) & (sk[88]) & (!g105)));
	assign g583 = (((!sk[89]) & (!g584) & (g585)) + ((sk[89]) & (!g584) & (!g585)));
	assign g584 = (((!sk[90]) & (!g359) & (g586)) + ((!sk[90]) & (!g359) & (g586)));
	assign g585 = (((!sk[91]) & (!g359) & (g589)) + ((!sk[91]) & (g359) & (g589)));
	assign g586 = (((!g587) & (!sk[92]) & (g588)) + ((!g587) & (sk[92]) & (!g588)));
	assign g587 = (((!i_6_) & (!sk[93]) & (g592)) + ((!i_6_) & (!sk[93]) & (g592)));
	assign g588 = (((!sk[94]) & (!i_6_) & (g593)) + ((!sk[94]) & (i_6_) & (g593)));
	assign g589 = (((!g590) & (!sk[95]) & (g591)) + ((!g590) & (sk[95]) & (!g591)));
	assign g590 = (((!i_6_) & (!sk[96]) & (g594)) + ((!i_6_) & (!sk[96]) & (g594)));
	assign g591 = (((i_6_) & (!sk[97]) & (g595)) + ((!i_6_) & (!sk[97]) & (g595)));
	assign g592 = (((!sk[98]) & (!i_8_) & (i_7_) & (!g105) & (!g392)) + ((!sk[98]) & (!i_8_) & (!i_7_) & (g105) & (!g392)) + ((!sk[98]) & (!i_8_) & (!i_7_) & (g105) & (g392)) + ((sk[98]) & (!i_8_) & (!i_7_) & (!g105) & (g392)) + ((!sk[98]) & (i_8_) & (i_7_) & (!g105) & (g392)));
	assign g593 = (((!sk[99]) & (!i_8_) & (i_7_) & (!g98) & (!g392)) + ((!sk[99]) & (!i_8_) & (!i_7_) & (g98) & (!g392)) + ((sk[99]) & (!i_8_) & (!i_7_) & (!g98) & (g392)) + ((!sk[99]) & (i_8_) & (!i_7_) & (g98) & (g392)));
	assign g594 = (((i_8_) & (!i_7_) & (!sk[100]) & (g392)) + ((!i_8_) & (!i_7_) & (!sk[100]) & (g392)) + ((!i_8_) & (!i_7_) & (!sk[100]) & (g392)));
	assign g595 = (((!i_8_) & (i_7_) & (!sk[101]) & (!g98) & (!g392)) + ((!i_8_) & (!i_7_) & (!sk[101]) & (g98) & (!g392)) + ((!i_8_) & (!i_7_) & (sk[101]) & (!g98) & (g392)) + ((i_8_) & (!i_7_) & (!sk[101]) & (g98) & (g392)));
	assign g596 = (((!sk[102]) & (!g597) & (g598)) + ((sk[102]) & (!g597) & (!g598)));
	assign g597 = (((!i_6_) & (!sk[103]) & (g599)) + ((!i_6_) & (!sk[103]) & (g599)));
	assign g598 = (((i_6_) & (!sk[104]) & (g601)) + ((!i_6_) & (!sk[104]) & (g601)));
	assign g599 = (((!i_7_) & (!sk[105]) & (g600)) + ((!i_7_) & (sk[105]) & (!g600)));
	assign g600 = (((!i_7_) & (!sk[106]) & (g604)) + ((!i_7_) & (!sk[106]) & (g604)));
	assign g601 = (((!sk[107]) & (!g602) & (g603)) + ((sk[107]) & (!g602) & (!g603)));
	assign g602 = (((!sk[108]) & (!i_7_) & (g605)) + ((!sk[108]) & (!i_7_) & (g605)));
	assign g603 = (((!sk[109]) & (!i_7_) & (g606)) + ((!sk[109]) & (i_7_) & (g606)));
	assign g604 = (((!g59) & (!sk[110]) & (!g25) & (i_8_)) + ((!g59) & (sk[110]) & (!g25) & (!i_8_)) + ((g59) & (!sk[110]) & (!g25) & (i_8_)) + ((!g59) & (!sk[110]) & (g25) & (i_8_)));
	assign g605 = (((!sk[111]) & (!g98) & (i_8_)) + ((sk[111]) & (!g98) & (!i_8_)) + ((!sk[111]) & (!g98) & (i_8_)));
	assign g606 = (((!sk[112]) & (!g25) & (g21)) + ((sk[112]) & (g25) & (!g21)));
	assign g607 = (((!sk[113]) & (!g608) & (g609)) + ((sk[113]) & (!g608) & (!g609)));
	assign g608 = (((!g6) & (!sk[114]) & (g610)) + ((!g6) & (!sk[114]) & (g610)));
	assign g609 = (((!sk[115]) & (!g6) & (g612)) + ((!sk[115]) & (g6) & (g612)));
	assign g610 = (((!sk[116]) & (!g11) & (g611)) + ((sk[116]) & (!g11) & (!g611)));
	assign g611 = (((!g11) & (!sk[117]) & (g615)) + ((!g11) & (!sk[117]) & (g615)));
	assign g612 = (((!g613) & (!sk[118]) & (g614)) + ((!g613) & (sk[118]) & (!g614)));
	assign g613 = (((!g11) & (!sk[119]) & (g616)) + ((!g11) & (!sk[119]) & (g616)));
	assign g614 = (((!sk[120]) & (!g11) & (g617)) + ((!sk[120]) & (g11) & (g617)));
	assign g615 = (((!sk[121]) & (!g13) & (g47)) + ((sk[121]) & (!g13) & (!g47)) + ((!sk[121]) & (g13) & (g47)));
	assign g616 = (((!g13) & (!sk[122]) & (g24) & (!g47) & (!g99)) + ((!g13) & (!sk[122]) & (!g24) & (g47) & (!g99)) + ((g13) & (!sk[122]) & (g24) & (!g47) & (!g99)) + ((!g13) & (!sk[122]) & (g24) & (!g47) & (!g99)));
	assign g617 = (((!g24) & (!g36) & (!sk[123]) & (g99)) + ((g24) & (!g36) & (sk[123]) & (!g99)) + ((!g24) & (g36) & (sk[123]) & (!g99)));
	assign g618 = (((!g619) & (!sk[124]) & (g620)) + ((!g619) & (sk[124]) & (!g620)));
	assign g619 = (((!g11) & (!sk[125]) & (g621)) + ((!g11) & (!sk[125]) & (g621)));
	assign g620 = (((g11) & (!sk[126]) & (g624)) + ((!g11) & (!sk[126]) & (g624)));
	assign g621 = (((!sk[127]) & (!g622) & (g623)) + ((sk[127]) & (!g622) & (!g623)));
	assign g622 = (((!sk[0]) & (!i_8_) & (g627)) + ((!sk[0]) & (!i_8_) & (g627)));
	assign g623 = (((!sk[1]) & (!i_8_) & (g628)) + ((!sk[1]) & (i_8_) & (g628)));
	assign g624 = (((!g625) & (!sk[2]) & (g626)) + ((!g625) & (sk[2]) & (!g626)));
	assign g625 = (((!sk[3]) & (!i_8_) & (g629)) + ((!sk[3]) & (!i_8_) & (g629)));
	assign g626 = (((!sk[4]) & (!i_8_) & (g630)) + ((!sk[4]) & (i_8_) & (g630)));
	assign g627 = (((!sk[5]) & (!i_6_) & (g46)) + ((sk[5]) & (!i_6_) & (!g46)) + ((!sk[5]) & (!i_6_) & (g46)));
	assign g628 = (((!g77) & (!i_6_) & (!sk[6]) & (i_7_) & (!g1)) + ((!g77) & (i_6_) & (!sk[6]) & (!i_7_) & (!g1)) + ((!g77) & (i_6_) & (!sk[6]) & (!i_7_) & (g1)) + ((!g77) & (!i_6_) & (sk[6]) & (!i_7_) & (!g1)));
	assign g629 = (((!sk[7]) & (!i_6_) & (g46)) + ((sk[7]) & (!i_6_) & (!g46)) + ((!sk[7]) & (!i_6_) & (g46)));
	assign g630 = (((!sk[8]) & (!g77) & (!i_6_) & (i_7_)) + ((sk[8]) & (!g77) & (!i_6_) & (!i_7_)) + ((sk[8]) & (!g77) & (i_6_) & (!i_7_)));
	assign g631 = (((!g632) & (!sk[9]) & (g633)) + ((!g632) & (sk[9]) & (!g633)));
	assign g632 = (((!sk[10]) & (!g35) & (g634)) + ((!sk[10]) & (!g35) & (g634)));
	assign g633 = (((!sk[11]) & (!g35) & (g637)) + ((!sk[11]) & (g35) & (g637)));
	assign g634 = (((!g635) & (!sk[12]) & (g636)) + ((!g635) & (sk[12]) & (!g636)));
	assign g635 = (((!i_5_) & (!sk[13]) & (g640)) + ((!i_5_) & (!sk[13]) & (g640)));
	assign g636 = (((!sk[14]) & (!i_5_) & (g641)) + ((!sk[14]) & (i_5_) & (g641)));
	assign g637 = (((!sk[15]) & (!g638) & (g639)) + ((sk[15]) & (!g638) & (!g639)));
	assign g638 = (((!sk[16]) & (!i_5_) & (g642)) + ((!sk[16]) & (!i_5_) & (g642)));
	assign g639 = (((!sk[17]) & (!i_5_) & (g643)) + ((!sk[17]) & (i_5_) & (g643)));
	assign g640 = (((!i_4_) & (!sk[18]) & (g121)) + ((!i_4_) & (sk[18]) & (!g121)) + ((!i_4_) & (!sk[18]) & (g121)));
	assign g641 = (((!g95) & (!sk[19]) & (!i_4_) & (i_6_)) + ((!g95) & (sk[19]) & (!i_4_) & (!i_6_)) + ((!g95) & (sk[19]) & (!i_4_) & (!i_6_)));
	assign g642 = (((!i_4_) & (!sk[20]) & (g121)) + ((!i_4_) & (sk[20]) & (!g121)) + ((!i_4_) & (!sk[20]) & (g121)));
	assign g643 = (((!g95) & (i_4_) & (!sk[21]) & (!i_6_) & (!g42)) + ((!g95) & (i_4_) & (!sk[21]) & (!i_6_) & (!g42)) + ((!g95) & (i_4_) & (!sk[21]) & (i_6_) & (!g42)) + ((!g95) & (!i_4_) & (!sk[21]) & (i_6_) & (!g42)) + ((!g95) & (!i_4_) & (sk[21]) & (!i_6_) & (!g42)));
	assign g644 = (((!g645) & (!sk[22]) & (g646)) + ((!g645) & (sk[22]) & (!g646)));
	assign g645 = (((!g42) & (!sk[23]) & (g647)) + ((!g42) & (!sk[23]) & (g647)));
	assign g646 = (((g42) & (!sk[24]) & (g650)) + ((!g42) & (!sk[24]) & (g650)));
	assign g647 = (((!g648) & (!sk[25]) & (g649)) + ((!g648) & (sk[25]) & (!g649)));
	assign g648 = (((!i_6_) & (!sk[26]) & (g653)) + ((!i_6_) & (!sk[26]) & (g653)));
	assign g649 = (((!sk[27]) & (!i_6_) & (g654)) + ((!sk[27]) & (i_6_) & (g654)));
	assign g650 = (((!sk[28]) & (!g651) & (g652)) + ((sk[28]) & (!g651) & (!g652)));
	assign g651 = (((!sk[29]) & (!i_6_) & (g655)) + ((!sk[29]) & (!i_6_) & (g655)));
	assign g652 = (((!sk[30]) & (!i_6_) & (g656)) + ((!sk[30]) & (i_6_) & (g656)));
	assign g653 = (((!g24) & (i_8_) & (!g36) & (!sk[31]) & (!i_7_)) + ((!g24) & (!i_8_) & (g36) & (!sk[31]) & (!i_7_)) + ((g24) & (!i_8_) & (!g36) & (sk[31]) & (!i_7_)) + ((!g24) & (!i_8_) & (!g36) & (sk[31]) & (i_7_)));
	assign g654 = (((!g24) & (!sk[32]) & (!i_8_) & (g45) & (!i_7_)) + ((!g24) & (!sk[32]) & (i_8_) & (!g45) & (!i_7_)) + ((!g24) & (sk[32]) & (!i_8_) & (!g45) & (!i_7_)) + ((g24) & (!sk[32]) & (i_8_) & (!g45) & (!i_7_)) + ((!g24) & (!sk[32]) & (i_8_) & (!g45) & (i_7_)));
	assign g655 = (((!sk[33]) & (!g24) & (i_8_) & (!g36) & (!i_7_)) + ((!sk[33]) & (!g24) & (!i_8_) & (g36) & (!i_7_)) + ((sk[33]) & (g24) & (!i_8_) & (!g36) & (!i_7_)) + ((sk[33]) & (!g24) & (!i_8_) & (!g36) & (i_7_)));
	assign g656 = (((!sk[34]) & (!g24) & (!i_8_) & (g45) & (!i_7_)) + ((!sk[34]) & (!g24) & (i_8_) & (!g45) & (!i_7_)) + ((!sk[34]) & (g24) & (i_8_) & (!g45) & (!i_7_)) + ((sk[34]) & (!g24) & (!i_8_) & (!g45) & (i_7_)));
	assign g657 = (((!g658) & (!sk[35]) & (g659)) + ((!g658) & (sk[35]) & (!g659)));
	assign g658 = (((!g23) & (!sk[36]) & (g660)) + ((!g23) & (!sk[36]) & (g660)));
	assign g659 = (((!sk[37]) & (!g23) & (g663)) + ((!sk[37]) & (g23) & (g663)));
	assign g660 = (((!g661) & (!sk[38]) & (g662)) + ((!g661) & (sk[38]) & (!g662)));
	assign g661 = (((!sk[39]) & (!i_2_) & (g666)) + ((!sk[39]) & (!i_2_) & (g666)));
	assign g662 = (((i_2_) & (!sk[40]) & (g667)) + ((!i_2_) & (!sk[40]) & (g667)));
	assign g663 = (((!g664) & (!sk[41]) & (g665)) + ((!g664) & (sk[41]) & (!g665)));
	assign g664 = (((!sk[42]) & (!i_2_) & (g668)) + ((!sk[42]) & (!i_2_) & (g668)));
	assign g665 = (((!sk[43]) & (!i_2_) & (g669)) + ((!sk[43]) & (i_2_) & (g669)));
	assign g666 = (((!i_0_) & (!g187) & (!sk[44]) & (i_1_) & (!g38)) + ((!i_0_) & (!g187) & (sk[44]) & (!i_1_) & (!g38)) + ((!i_0_) & (g187) & (!sk[44]) & (!i_1_) & (!g38)) + ((!i_0_) & (g187) & (!sk[44]) & (!i_1_) & (g38)));
	assign g667 = (((!i_0_) & (!i_7_) & (!sk[45]) & (g38)) + ((!i_0_) & (!i_7_) & (sk[45]) & (!g38)) + ((!i_0_) & (!i_7_) & (sk[45]) & (!g38)));
	assign g668 = (((!i_0_) & (!g187) & (!sk[46]) & (i_1_)) + ((!i_0_) & (!g187) & (sk[46]) & (!i_1_)) + ((!i_0_) & (g187) & (sk[46]) & (!i_1_)));
	assign g669 = (((!sk[47]) & (!i_0_) & (!i_7_) & (g38)) + ((sk[47]) & (!i_0_) & (!i_7_) & (!g38)) + ((sk[47]) & (!i_0_) & (!i_7_) & (!g38)));
	assign g670 = (((!sk[48]) & (!g671) & (g672)) + ((sk[48]) & (!g671) & (!g672)));
	assign g671 = (((!sk[49]) & (!g41) & (g673)) + ((!sk[49]) & (!g41) & (g673)));
	assign g672 = (((g41) & (!sk[50]) & (g676)) + ((!g41) & (!sk[50]) & (g676)));
	assign g673 = (((!g674) & (!sk[51]) & (g675)) + ((!g674) & (sk[51]) & (!g675)));
	assign g674 = (((!i_4_) & (!sk[52]) & (g679)) + ((!i_4_) & (!sk[52]) & (g679)));
	assign g675 = (((!sk[53]) & (!i_4_) & (g680)) + ((!sk[53]) & (i_4_) & (g680)));
	assign g676 = (((!g677) & (!sk[54]) & (g678)) + ((!g677) & (sk[54]) & (!g678)));
	assign g677 = (((!i_4_) & (!sk[55]) & (g681)) + ((!i_4_) & (!sk[55]) & (g681)));
	assign g678 = (((i_4_) & (!sk[56]) & (g682)) + ((!i_4_) & (!sk[56]) & (g682)));
	assign g679 = (((!g1) & (i_5_) & (!g12) & (!sk[57]) & (!i_3_)) + ((!g1) & (!i_5_) & (!g12) & (sk[57]) & (!i_3_)) + ((!g1) & (!i_5_) & (g12) & (!sk[57]) & (!i_3_)) + ((g1) & (!i_5_) & (!g12) & (sk[57]) & (!i_3_)) + ((!g1) & (!i_5_) & (!g12) & (sk[57]) & (!i_3_)));
	assign g680 = (((!g1) & (!sk[58]) & (i_5_) & (!g28) & (!i_3_)) + ((!g1) & (!sk[58]) & (!i_5_) & (g28) & (!i_3_)) + ((!g1) & (sk[58]) & (!i_5_) & (!g28) & (!i_3_)) + ((g1) & (!sk[58]) & (!i_5_) & (g28) & (!i_3_)) + ((!g1) & (!sk[58]) & (!i_5_) & (g28) & (!i_3_)));
	assign g681 = (((!g1) & (i_5_) & (!sk[59]) & (!g12) & (!i_3_)) + ((!g1) & (!i_5_) & (!sk[59]) & (g12) & (!i_3_)) + ((!g1) & (!i_5_) & (sk[59]) & (!g12) & (i_3_)) + ((g1) & (!i_5_) & (!sk[59]) & (g12) & (i_3_)));
	assign g682 = (((!sk[60]) & (!g1) & (i_5_) & (!g28) & (!i_3_)) + ((!sk[60]) & (!g1) & (!i_5_) & (g28) & (!i_3_)) + ((sk[60]) & (!g1) & (!i_5_) & (!g28) & (!i_3_)) + ((!sk[60]) & (g1) & (!i_5_) & (g28) & (!i_3_)) + ((!sk[60]) & (!g1) & (!i_5_) & (g28) & (!i_3_)));
	assign g683 = (((!sk[61]) & (!g684) & (g685)) + ((sk[61]) & (!g684) & (!g685)));
	assign g684 = (((!g27) & (!sk[62]) & (g686)) + ((!g27) & (!sk[62]) & (g686)));
	assign g685 = (((g27) & (!sk[63]) & (g689)) + ((!g27) & (!sk[63]) & (g689)));
	assign g686 = (((!g687) & (!sk[64]) & (g688)) + ((!g687) & (sk[64]) & (!g688)));
	assign g687 = (((!i_8_) & (!sk[65]) & (g691)) + ((!i_8_) & (!sk[65]) & (g691)));
	assign g688 = (((i_8_) & (!sk[66]) & (g692)) + ((!i_8_) & (!sk[66]) & (g692)));
	assign g689 = (((!i_8_) & (!sk[67]) & (g690)) + ((!i_8_) & (sk[67]) & (!g690)));
	assign g690 = (((!i_8_) & (!sk[68]) & (g693)) + ((!i_8_) & (!sk[68]) & (g693)));
	assign g691 = (((!g116) & (i_7_) & (!sk[69]) & (!g126) & (!i_6_)) + ((!g116) & (!i_7_) & (!sk[69]) & (g126) & (!i_6_)) + ((!g116) & (!i_7_) & (!sk[69]) & (g126) & (i_6_)) + ((!g116) & (!i_7_) & (sk[69]) & (!g126) & (!i_6_)));
	assign g692 = (((!g116) & (!i_7_) & (g5) & (!sk[70]) & (!i_6_)) + ((!g116) & (i_7_) & (!g5) & (!sk[70]) & (!i_6_)) + ((!g116) & (i_7_) & (!g5) & (!sk[70]) & (!i_6_)) + ((!g116) & (!i_7_) & (!g5) & (sk[70]) & (!i_6_)) + ((!g116) & (!i_7_) & (!g5) & (sk[70]) & (i_6_)));
	assign g693 = (((!i_7_) & (!g126) & (!sk[71]) & (i_6_)) + ((!i_7_) & (!g126) & (sk[71]) & (!i_6_)) + ((i_7_) & (!g126) & (!sk[71]) & (i_6_)) + ((!i_7_) & (g126) & (!sk[71]) & (i_6_)));
	assign g694 = (((!sk[72]) & (!g695) & (g696)) + ((sk[72]) & (!g695) & (!g696)));
	assign g695 = (((!g47) & (!sk[73]) & (g697)) + ((!g47) & (!sk[73]) & (g697)));
	assign g696 = (((g47) & (!sk[74]) & (g699)) + ((!g47) & (!sk[74]) & (g699)));
	assign g697 = (((!sk[75]) & (!i_4_) & (g698)) + ((sk[75]) & (!i_4_) & (!g698)));
	assign g698 = (((!sk[76]) & (!i_4_) & (g702)) + ((!sk[76]) & (!i_4_) & (g702)));
	assign g699 = (((!g700) & (!sk[77]) & (g701)) + ((!g700) & (sk[77]) & (!g701)));
	assign g700 = (((!sk[78]) & (!i_4_) & (g703)) + ((!sk[78]) & (!i_4_) & (g703)));
	assign g701 = (((!sk[79]) & (!i_4_) & (g704)) + ((!sk[79]) & (i_4_) & (g704)));
	assign g702 = (((!i_5_) & (!sk[80]) & (!g121) & (i_3_)) + ((!i_5_) & (sk[80]) & (!g121) & (!i_3_)) + ((!i_5_) & (sk[80]) & (!g121) & (!i_3_)));
	assign g703 = (((!i_5_) & (!sk[81]) & (!g121) & (i_3_)) + ((!i_5_) & (sk[81]) & (!g121) & (!i_3_)) + ((!i_5_) & (sk[81]) & (!g121) & (!i_3_)));
	assign g704 = (((!i_6_) & (!sk[82]) & (!i_5_) & (g27) & (!i_3_)) + ((!i_6_) & (!sk[82]) & (i_5_) & (!g27) & (!i_3_)) + ((!i_6_) & (!sk[82]) & (i_5_) & (!g27) & (!i_3_)) + ((!i_6_) & (sk[82]) & (!i_5_) & (!g27) & (!i_3_)) + ((i_6_) & (sk[82]) & (!i_5_) & (!g27) & (!i_3_)));
	//assign gnd = ();

endmodule