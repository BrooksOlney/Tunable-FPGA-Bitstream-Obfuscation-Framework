module s38417 (
	Pg3234, Pg3233, Pg3232, Pg3231, Pg3230, Pg3229, Pg3228, Pg3227, 
	Pg3226, Pg3225, Pg3224, Pg3223, Pg3222, Pg3221, Pg3220, Pg3219, Pg3218, Pg3217, 
	Pg3216, Pg3215, Pg3214, Pg3213, Pg3212, Pg2637, Pg1943, Pg1249, Pg563, Pg51, 
	PCLK, Pg27380, Pg26149, Pg26135, Pg26104, Pg25489, Pg25442, Pg25435, Pg25420, Pg24734, 
	Pg16496, Pg16437, Pg16399, Pg16355, Pg16297, Pg8275, Pg8274, Pg8273, Pg8272, Pg8271, 
	Pg8270, Pg8269, Pg8268, Pg8267, Pg8266, Pg8265, Pg8264, Pg8263, Pg8262, Pg8261, 
	Pg8260, Pg8259, Pg8258, Pg8251, Pg8249, Pg8175, Pg8167, Pg8106, Pg8096, Pg8087, 
	Pg8082, Pg8030, Pg8023, Pg8021, Pg8012, Pg8007, Pg7961, Pg7956, Pg7909, Pg7519, 
	Pg7487, Pg7425, Pg7390, Pg7357, Pg7334, Pg7302, Pg7264, Pg7229, Pg7194, Pg7161, 
	Pg7084, Pg7052, Pg7014, Pg6979, Pg6944, Pg6911, Pg6895, Pg6837, Pg6782, Pg6750, 
	Pg6712, Pg6677, Pg6642, Pg6573, Pg6518, Pg6485, Pg6447, Pg6442, Pg6368, Pg6313, 
	Pg6231, Pg6225, Pg5796, Pg5747, Pg5738, Pg5695, Pg5686, Pg5657, Pg5648, Pg5637, 
	Pg5629, Pg5612, Pg5595, Pg5555, Pg5549, Pg5511, Pg5472, Pg5437, Pg5388, Pg4590, 
	Pg4450, Pg4323, Pg4321, Pg4200, Pg4090, Pg4088, Pg3993);

input Pg3234, Pg3233, Pg3232, Pg3231, Pg3230, Pg3229, Pg3228, Pg3227, Pg3226, Pg3225, Pg3224, Pg3223, Pg3222, Pg3221, Pg3220, Pg3219, Pg3218, Pg3217, Pg3216, Pg3215, Pg3214, Pg3213, Pg3212, Pg2637, Pg1943, Pg1249, Pg563, Pg51, PCLK;

output Pg27380, Pg26149, Pg26135, Pg26104, Pg25489, Pg25442, Pg25435, Pg25420, Pg24734, Pg16496, Pg16437, Pg16399, Pg16355, Pg16297, Pg8275, Pg8274, Pg8273, Pg8272, Pg8271, Pg8270, Pg8269, Pg8268, Pg8267, Pg8266, Pg8265, Pg8264, Pg8263, Pg8262, Pg8261, Pg8260, Pg8259, Pg8258, Pg8251, Pg8249, Pg8175, Pg8167, Pg8106, Pg8096, Pg8087, Pg8082, Pg8030, Pg8023, Pg8021, Pg8012, Pg8007, Pg7961, Pg7956, Pg7909, Pg7519, Pg7487, Pg7425, Pg7390, Pg7357, Pg7334, Pg7302, Pg7264, Pg7229, Pg7194, Pg7161, Pg7084, Pg7052, Pg7014, Pg6979, Pg6944, Pg6911, Pg6895, Pg6837, Pg6782, Pg6750, Pg6712, Pg6677, Pg6642, Pg6573, Pg6518, Pg6485, Pg6447, Pg6442, Pg6368, Pg6313, Pg6231, Pg6225, Pg5796, Pg5747, Pg5738, Pg5695, Pg5686, Pg5657, Pg5648, Pg5637, Pg5629, Pg5612, Pg5595, Pg5555, Pg5549, Pg5511, Pg5472, Pg5437, Pg5388, Pg4590, Pg4450, Pg4323, Pg4321, Pg4200, Pg4090, Pg4088, Pg3993;

wire wire1521, n1139, n1138, n1137, n1142, n1141, n1140, n1145, n1144, n1143, n1148, n1147, n1146, n69, n66, n72, n70, n75, n73, n78, n76, n81, n79, n84, n82, n87, n85, n90, n88, n93, n91, n96, n94, n99, n97, n102, n100, n105, n103, n108, n106, n111, n109, n114, n112, n117, n115, n120, n118, n123, n121, n126, n124, n129, n127, n131, n130, n133, Ng19021, n134, Ng19022, n136, n135, n138, n137, n139, Ng19033, n140, Ng19023, n141, Ng19034, n143, n142, n145, n144, n146, Ng19045, n148, Ng16467, n149, Ng19035, n150, Ng19046, n152, n151, n154, n153, n155, Ng19057, n157, Ng16469, n158, Ng19047, n159, Ng19058, n161, n160, n163, Ng16471, n164, Ng19059, n166, Ng16468, n168, n167, n170, Ng16473, n172, Ng16470, n174, n173, n176, Ng16472, n178, n177, n180, Ng16474, n183, n181, n185, n184, n187, n186, n188, n190, n189, n192, n191, n194, n193, n196, n195, n199, n197, n201, n200, n203, n202, n205, n204, n207, n206, n211, n208, n213, n212, n216, n214, n218, n217, n220, n219, n222, n221, n225, n223, n227, n226, n229, n228, n231, n230, n234, n232, n236, n235, n239, n237, n241, n240, n243, n242, n246, n244, n248, n247, n250, n249, n253, n251, n255, n254, n257, n256, n259, n258, n262, n260, n264, n263, n267, n265, n269, n268, n271, n270, n274, n272, n276, n275, n278, n277, n281, n279, n283, n282, n285, n284, n288, n286, n290, n289, n292, n291, n294, n293, n297, n295, n299, n298, n302, n300, n304, n303, n307, n305, n309, n308, n311, n310, n313, n312, n316, n314, n318, n317, n320, n319, n323, n321, n325, n324, n327, n326, n330, n328, n332, n331, n334, n333, n337, n335, n340, n338, n342, n341, n345, n343, n347, n346, n349, n348, n352, n350, n354, n353, n357, n355, n359, n358, n361, n360, n363, n362, n366, n364, n368, n367, n370, n369, n373, n371, n375, n374, n378, n376, n380, n379, n382, n381, n384, n383, n387, n385, n390, n388, n392, n391, n395, n393, n397, n396, n399, n398, n402, n400, n404, n403, n407, n405, n409, n408, n411, n410, n413, n412, n416, n414, n418, n417, n421, n419, n423, n422, n425, n424, n428, n426, n430, n429, n432, n431, n434, n433, n437, n435, n440, n438, n442, n441, n445, n443, n447, n446, n449, n448, n452, n450, n454, n453, n457, n455, n459, n458, n461, n460, n463, n462, n466, n464, n468, n467, n470, n469, n473, n471, n475, n474, n477, n476, n479, n478, n482, n480, n485, n483, n487, n486, n490, n488, n492, n491, n494, n493, n496, n495, n498, n497, n501, n499, n503, n502, n505, n504, n508, n506, n510, n509, n512, n511, n514, n513, n516, n515, n518, n517, n520, n519, n523, n521, n525, n524, n527, n526, n529, n528, n531, n530, n533, n532, n535, n534, n537, n536, n539, n538, n541, n540, n543, n542, n545, n544, n547, n546, n550, n548, n552, n551, n554, n553, n556, n555, n559, n557, n561, n560, n563, n562, n566, n564, n568, n567, n571, n569, n573, n572, n575, n574, n577, n576, n580, n578, n582, n581, n584, n583, n586, n585, n589, n587, n591, n590, n594, n592, n596, n595, n598, n597, n600, n599, n603, n601, n605, n604, n608, n606, n610, n609, n612, n611, n614, n613, n617, n615, n619, n618, n622, n620, n624, n623, n626, n625, n628, n627, n631, n629, n633, n632, n635, n634, n637, n636, n639, n638, n641, n640, n643, n642, n644, Ng16494, n646, n645, n648, n647, n651, n649, n653, n652, n656, n654, n658, n657, n661, n659, n664, n662, n665, n667, n669, n671, n673, n675, n677, n679, n683, n684, n681, n687, n688, n685, n691, n692, n689, n695, n696, n693, Ng20571, Ng20588, n698, Ng21943, n699, Ng21944, n700, Ng21945, n701, Ng21946, Ng21951, Ng21965, n702, Ng23160, n703, Ng23198, n704, Ng23236, n705, Ng23274, n706, n707, Ng23161, n708, n709, Ng23199, n710, n711, Ng23237, n712, n713, Ng23275, n714, n715, Ng23315, Ng23317, Ng23318, n717, Ng24296, n718, Ng24337, n722, n721, n719, n723, Ng24378, n726, n724, n727, Ng24419, n730, n728, n733, n731, n734, n735, Ng24424, n736, Ng24295, n737, n738, Ng24425, n739, Ng24336, n740, Ng24377, n742, Ng24423, n744, n743, Ng24297, n745, Ng24418, n746, Ng24298, n748, n747, Ng24338, n750, n749, n752, n751, Ng24299, n753, Ng24339, n755, n754, Ng24379, n757, n756, n759, n758, Ng24340, n760, Ng24380, n762, n761, Ng24420, n764, n763, n766, n765, Ng24381, n767, Ng24421, n769, n768, n771, n770, Ng24422, Ng28313, n772, Ng25140, n773, Ng25151, n775, Ng25177, n776, Ng25162, n777, Ng25173, n778, Ng25174, n780, Ng25175, n781, Ng25176, Ng28696, n783, Ng25991, n784, Ng26000, n785, Ng26009, n786, Ng26018, n787, Ng26021, n788, Ng26022, n789, Ng26019, n790, Ng26020, n791, n792, Ng26678, n793, Ng26695, n794, Ng26712, n795, Ng26729, Ng29166, n796, Ng26691, n797, Ng26708, n798, Ng26750, n799, Ng26725, n800, Ng26742, n801, Ng26746, n802, Ng26747, n803, Ng26749, n804, Ng27189, n805, Ng27198, n806, Ng27219, n807, Ng27228, n808, Ng27197, n809, Ng27218, n810, Ng27227, n811, Ng27236, n812, Ng27239, n813, Ng27237, n814, Ng27683, n815, Ng27691, n816, Ng27699, n817, Ng27707, Ng29656, n818, Ng27690, n819, Ng27698, Ng27716, n821, Ng27706, n822, Ng27714, n823, Ng27715, n824, Ng28206, n825, Ng28232, n826, Ng28258, n827, Ng28284, n828, Ng28231, n829, Ng28257, n830, Ng28283, n831, Ng28309, n833, n834, n832, n836, n837, n835, n839, n840, n838, n842, n843, n841, n844, Ng28673, n845, Ng28678, n846, Ng28683, n847, Ng28688, n848, Ng28677, n849, Ng28682, n850, Ng28687, n851, Ng28692, n852, n853, Ng28674, n854, Ng28675, n855, n856, Ng28679, n857, Ng28676, n858, Ng28680, n859, n860, Ng28684, n861, Ng28681, n862, Ng28685, n863, n864, Ng28689, n865, Ng28686, n866, Ng28690, n867, Ng28691, n868, Ng29131, n869, Ng29139, n870, Ng29147, n871, Ng29155, n872, Ng29138, n873, Ng29146, n874, Ng29154, n875, Ng29162, n876, Ng29413, n877, Ng29420, n878, Ng29427, n879, Ng29446, n881, n880, Ng29417, n882, Ng29418, n884, n883, Ng29424, n885, Ng29419, n886, Ng29425, n888, n887, Ng29437, n889, Ng29426, n890, Ng29438, n892, n891, Ng29450, n893, Ng29439, n894, Ng29451, n895, Ng29452, n896, Ng29627, n897, Ng29634, n898, Ng29641, n899, Ng29648, n900, Ng29794, n901, Ng29798, n902, Ng29802, n903, Ng29806, n907, n908, n904, n912, n913, n909, n917, n918, n914, n922, n923, n919, n925, n927, n924, n930, n931, n929, n933, n935, n932, n938, n939, n937, n941, n942, n940, n944, n946, n943, n949, n950, n948, n952, n953, n951, n955, n957, n954, n960, n961, n959, n963, n964, n962, n966, n967, n965, n969, n970, n968, n972, n973, n971, n975, n976, n974, n978, n979, n977, n981, n982, n980, n984, n985, n983, n987, n988, n986, n990, n991, n989, n994, n993, n992, n997, n996, n1000, n999, n1004, n1002, n1005, n1008, n1007, n1010, n1009, n1012, n1011, n1015, n1013, n1019, n1017, n1023, n1022, n1021, n1025, n1024, n1028, n1027, n1031, n1030, n1032, n1035, n1034, n1037, n1036, n1039, n1038, n1043, n1042, n1047, n1046, n1051, n1050, n1056, n1054, n1059, n1058, n1062, n1061, n1065, n1064, n1068, n1067, n1072, n1070, n1074, n1073, n1076, n1075, n1078, n1077, n1081, n1080, n1084, n1083, n1085, n1088, n1087, n1091, n1089, n1094, n1093, n1098, n1096, n1100, n1099, n1102, n1101, n1104, n1103, n1107, n1106, n1110, n1109, n1111, n1115, n1113, n1118, n1119, n1120, n1121, n1117, n1123, n1124, n1125, n1126, n1122, n1128, n1129, n1130, n1131, n1127, n1133, n1134, n1135, n1136, n1132, n1149, n1151, n1154, n1155, n1156, n1157, n1153, n1159, n1160, n1161, n1162, n1158, n1163, n1165, n1168, n1169, n1170, n1171, n1167, n1173, n1174, n1175, n1176, n1172, n1177, n1179, n1182, n1183, n1184, n1185, n1181, n1187, n1188, n1189, n1190, n1186, n1191, n1193, n1196, n1197, n1198, n1199, n1195, n1201, n1202, n1203, n1204, n1200, n1207, n1206, n1205, n1210, n1209, n1208, n1213, n1212, n1211, n1216, n1215, n1214, Ng19048, Ng19036, Ng19024, Ng19012, n1217, Ng30989, n1218, Ng30987, n1219, Ng30986, n1220, Ng30985, n1221, Ng30984, n1222, Ng30983, n1223, Ng30982, n1224, Ng30981, n1225, Ng30980, n1226, Ng30940, n1227, Ng30915, n1228, Ng30914, n1229, Ng30913, n1230, Ng30912, n1231, Ng30911, n1232, Ng30910, n1233, Ng30909, n1234, Ng30908, n1235, Ng30119, n1236, Ng29979, n1237, Ng29978, n1238, Ng29977, n1239, Ng29976, n1240, Ng29975, n1241, Ng29974, n1242, Ng29973, n1243, Ng29972, n1244, Ng29655, n1245, Ng29460, n1246, Ng29459, n1247, Ng29458, n1248, Ng29457, n1249, Ng29456, n1250, Ng29455, n1251, Ng29454, n1252, Ng29453, Ng13466, Ng13465, Ng13464, Ng13463, Ng13462, Ng13461, Ng13460, Ng13459, Ng13458, Ng11576, Ng11575, Ng11574, Ng11573, Ng11572, Ng11592, Ng11591, Ng11590, Ng13450, Ng13449, Ng13448, Ng13447, Ng13446, Ng13445, Ng13444, Ng13443, Ng13442, Ng11549, Ng11548, Ng11547, Ng11546, Ng11545, Ng11565, Ng11564, Ng11563, Ng13434, Ng13433, Ng13432, Ng13431, Ng13430, Ng13429, Ng13428, Ng13427, Ng13426, Ng11522, Ng11521, Ng11520, Ng11519, Ng11518, Ng11538, Ng11537, Ng11536, Ng13418, Ng13417, Ng13416, Ng13415, Ng13414, Ng13413, Ng13412, Ng13411, Ng13410, Ng11495, Ng11494, Ng11493, Ng11492, Ng11491, Ng11511, Ng11510, Ng11509, n1254, n1253, n1256, n1257, n1255, n1259, n1260, n1258, n1262, n1263, n1261, n1264, n1267, n1270, n1273, n1282, n1276, n1284, n1283, n1287, n1290, n1293, n1306, n1300, n1308, n1307, n1311, n1314, n1316, n1324, n1325, n1323, n1329, n1330, n1328, n1333, n1334, n1332, n1339, n1338, n1340, n1341, n1343, n1344, n1342, n1345, n1349, n1352, n1351, n1357, n1358, n1356, n1362, n1363, n1361, n1366, n1367, n1365, n1372, n1371, n1373, n1374, n1376, n1377, n1375, n1378, n1382, n1385, n1384, n1390, n1391, n1389, n1395, n1396, n1394, n1399, n1400, n1398, n1405, n1404, n1406, n1407, n1409, n1410, n1408, n1411, n1415, n1418, n1417, n1423, n1424, n1422, n1428, n1429, n1427, n1432, n1433, n1431, n1438, n1437, n1439, n1440, n1442, n1443, n1441, n1444, n1448, n1451, n1450, n1457, n1455, n1458, n1459, n1460, n1461, n1462, n1465, n1463, n1466, n1467, n1468, n1469, n1470, n1473, n1471, n1474, n1475, n1476, n1477, n1478, n1481, n1479, n1482, n1483, n1484, n1485, n1486, n1488, n1487, n1491, n1490, n1494, n1497, n1500, n1507, n1510, n1509, n1511, n1514, n1513, n1515, n1518, n1517, n1519, n1522, n1521, n1526, n1524, n1525, n1523, n1529, n1527, n1530, n1533, n1532, n1536, n1535, n1541, n1538, n1539, n1540, n1537, n1545, n1546, n1542, n1551, n1548, n1549, n1550, n1547, n1555, n1556, n1552, n1561, n1558, n1559, n1560, n1557, n1565, n1566, n1562, n1571, n1568, n1569, n1570, n1567, n1575, n1576, n1572, n1579, n1582, n1585, n1595, n1593, n1598, n1597, n1602, n1600, n1605, n1604, n1609, n1607, n1612, n1611, n1616, n1614, n1619, n1618, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1629, n1628, n1630, n1634, n1636, n1640, n1639, n1641, n1646, n1644, n1647, n1648, n1650, n1653, n1654, n1652, n1657, n1658, n1656, n1661, n1662, n1659, n1664, n1663, n1665, n1669, n1671, n1675, n1674, n1676, n1681, n1679, n1682, n1683, n1685, n1688, n1689, n1687, n1692, n1693, n1691, n1696, n1697, n1694, n1699, n1698, n1700, n1704, n1706, n1710, n1709, n1711, n1716, n1714, n1717, n1718, n1720, n1723, n1724, n1722, n1727, n1728, n1726, n1731, n1732, n1729, n1734, n1733, n1735, n1739, n1741, n1745, n1744, n1746, n1751, n1749, n1752, n1753, n1755, n1758, n1759, n1757, n1762, n1763, n1761, n1766, n1767, n1764, n1768, n1769, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1770, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1778, n1789, n1786, n1791, n1792, n1790, n1796, n1795, n1800, n1797, n1802, n1803, n1801, n1806, n1805, n1810, n1807, n1812, n1813, n1811, n1816, n1815, n1820, n1817, n1822, n1823, n1821, n1826, n1825, n1830, n1834, n1831, n1837, n1835, n1840, n1843, n1841, n1846, n1844, n1849, n1852, n1850, n1855, n1853, n1858, n1861, n1859, n1864, n1862, n1867, n1865, n1869, n1868, n1871, n1870, n1873, n1872, n1875, n1874, n1877, n1876, n1879, n1878, n1881, n1880, n1883, n1882, n1885, n1884, n1886, n1887, n1889, Ng27229, n1890, n1891, n1893, Ng27220, n1894, n1895, n1897, Ng27199, n1898, n1899, n1901, Ng27190, n1902, n1905, n1907, n1906, n1908, n1912, n1911, n1914, n1913, n1916, n1915, n1919, n1918, n1920, n1923, n1922, n1924, n1927, n1926, n1928, n1930, n1934, n1933, n1936, n1935, n1938, n1937, n1940, n1939, n1942, n1941, n1944, n1943, n1946, n1945, n1947, n1948, n1951, n1949, n1952, n1954, n1956, n1960, n1958, n1966, n1968, n1970, n1972, n1976, n1974, n1978, Ng27238, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1998, n2000, n2002, n2003, n2005, n2006, n2008, n2009, n2011, n2012, n2014, n2015, n2017, n2018, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2031, n2033, n2035, n2036, n2038, n2039, n2041, n2042, n2044, n2045, n2047, n2048, n2050, n2051, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2064, n2066, n2068, n2069, n2071, n2072, n2074, n2075, n2077, n2078, n2080, n2081, n2083, n2084, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2097, n2099, n2101, n2102, n2104, n2105, n2107, n2108, n2110, n2111, n2113, n2114, n2116, n2117, n2119, n2121, n2120, n2123, n2122, n2125, n2124, n2127, n2126, n2138, n2139, n2140, n2141, n2143, n2142, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2189, n2191, n2192, n2194, n2196, n2198, n2199, n2201, n2203, n2204, n2205, n2207, n2208, n2210, n2212, n2214, n2215, n2217, n2219, n2220, n2221, n2223, n2225, n2227, n2229, n2231, n2233, n2235, n2237, n2239, n2241, n2243, n2245, n2247, n2249, n2251, n2253, n2255, n2257, n2259, Ng30325, n2278, Ng29445, n2291, n2295, n2296, n2297, n2319, n2320, n2323, n2324, n2325, n2326, n2327, n2330, n2331, n2332, n2354, n2355, n2358, n2359, n2360, n2361, n2362, n2365, n2366, n2367, n2389, n2390, n2393, n2394, n2395, n2396, n2397, n2400, n2401, n2402, n2424, n2425, n2428, n2429, n2430, n2431, n2432, Ng27217, n2444, n2450, n2453, n2455, n2460, Ng23159, n2467, n2489, n2491, n2493, n2495, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2508, n2510, n2512, n2514, n2515, n2517, n2519, n2520, n2521, n2523, n2524, n2534, n2546, n2545, n2547, n2551, n2560, n2572, n2571, n2575, n2584, n2596, n2595, n2599, n2608, n2620, n2619, n2653, n2662, n2671, n2680, n2694, n2695, n2699, n2702, n2703, n2704, n2705, n2706, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2721, Ng21966, n2722, Ng21964, Ng20604, Ng20594, n2724, Ng19061, n2725, Ng19060, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, Ng30943, n2736, Ng30942, n2737, Ng30941, n2738, n2739, n2740, n2741, n2742, n2743, Ng30907, n2744, Ng30906, n2745, Ng30905, n2746, n2747, n2748, Ng30904, n2749, Ng30903, n2750, Ng30902, n2751, Ng30901, n2752, Ng30900, n2753, Ng30899, n2754, Ng30898, n2755, Ng30897, n2756, Ng30896, n2757, Ng30895, n2758, Ng30894, n2759, Ng30893, n2760, Ng30892, n2761, Ng30891, n2762, Ng30890, n2763, Ng30889, n2764, Ng30888, n2765, Ng30887, n2766, n2767, n2768, Ng30886, n2769, Ng30885, n2770, Ng30884, n2771, Ng30883, n2772, Ng30882, n2773, Ng30881, n2774, Ng30880, n2775, Ng30879, n2776, Ng30878, n2777, Ng30877, n2778, Ng30876, n2779, Ng30875, n2780, Ng30874, n2781, Ng30873, n2782, Ng30872, n2783, Ng30871, n2784, Ng30870, n2785, Ng30869, n2786, n2787, n2788, Ng30868, n2789, Ng30867, n2790, Ng30866, n2791, Ng30865, n2792, Ng30864, n2793, Ng30863, n2794, Ng30862, n2795, Ng30861, n2796, Ng30860, n2797, Ng30859, n2798, Ng30858, n2799, Ng30857, n2800, Ng30856, n2801, Ng30855, n2802, Ng30854, n2803, Ng30853, n2804, Ng30852, n2805, Ng30851, n2806, n2807, n2808, Ng30850, n2809, Ng30849, n2810, Ng30848, n2811, Ng30847, n2812, Ng30846, n2813, Ng30845, n2814, Ng30844, n2815, Ng30843, n2816, Ng30842, n2817, Ng30841, n2818, Ng30840, n2819, Ng30839, n2820, Ng30838, n2821, Ng30837, n2822, Ng30836, n2823, Ng30721, n2824, Ng30720, n2825, Ng30719, n2826, Ng30718, n2827, Ng30717, n2828, Ng30716, n2829, Ng30715, n2830, Ng30714, n2831, Ng30713, n2832, Ng30712, n2833, Ng30711, n2834, Ng30710, n2836, n2837, Ng30565, n2838, Ng30564, n2839, Ng30563, n2840, Ng30562, n2841, Ng30561, n2842, Ng30560, n2844, n2845, Ng30559, n2846, Ng30558, n2847, Ng30557, n2849, n2850, Ng30556, n2851, Ng30555, n2852, Ng30554, n2854, n2855, Ng30553, n2856, Ng30552, n2857, Ng30551, n2859, n2860, Ng30550, n2861, Ng30549, n2862, Ng30548, n2863, Ng30547, n2864, Ng30546, n2865, Ng30545, n2867, n2868, Ng30544, n2869, Ng30543, n2870, Ng30542, n2872, n2873, Ng30541, n2874, Ng30540, n2875, Ng30539, n2877, n2878, Ng30538, n2879, Ng30537, n2880, Ng30536, n2882, n2883, Ng30535, n2884, Ng30534, n2885, Ng30533, n2886, Ng30532, n2887, Ng30531, n2888, Ng30530, n2890, n2891, Ng30529, n2892, Ng30528, n2893, Ng30527, n2895, n2896, Ng30526, n2897, Ng30525, n2898, Ng30524, n2900, n2901, Ng30523, n2902, Ng30522, n2903, Ng30521, n2905, n2906, Ng30520, n2907, Ng30519, n2908, Ng30518, n2909, Ng30517, n2910, Ng30516, n2911, Ng30515, n2913, n2914, Ng30514, n2915, Ng30513, n2916, Ng30512, n2918, n2919, Ng30511, n2920, Ng30510, n2921, Ng30509, n2923, n2924, Ng30508, n2925, Ng30507, n2926, Ng30506, Ng29440, n2928, Ng30320, n2929, Ng23148, n2930, Ng27200, n2931, Ng29428, n2932, Ng30314, n2933, Ng30122, n2934, Ng30121, n2935, Ng30120, n2936, n2937, n2938, n2939, n2940, n2941, Ng29809, n2942, Ng29808, n2943, Ng29807, n2944, Ng29805, n2945, Ng29804, n2946, Ng29803, n2947, Ng29801, n2948, Ng29800, n2949, Ng29799, n2950, Ng29797, n2951, Ng29796, n2952, Ng29795, n2954, n2955, n2956, n2957, n2958, n2959, n2960, Ng29654, n2961, Ng29653, n2962, Ng29652, n2963, Ng29651, n2964, Ng29650, n2965, Ng29649, n2966, Ng29647, n2967, Ng29646, n2968, Ng29645, n2969, Ng29644, n2970, Ng29643, n2971, Ng29642, n2972, Ng29640, n2973, Ng29639, n2974, Ng29638, n2975, Ng29637, n2976, Ng29636, n2977, Ng29635, n2978, Ng29633, n2979, Ng29632, n2980, Ng29631, n2981, Ng29630, n2982, Ng29629, n2983, Ng29628, n2984, Ng29449, n2985, Ng29448, n2986, Ng29447, n2987, Ng29436, n2988, Ng29435, n2989, Ng29434, n2990, Ng29423, n2991, Ng29422, n2992, Ng29421, n2993, Ng29416, n2994, Ng29415, n2995, Ng29414, n2996, Ng29165, n2997, Ng29164, n2998, Ng29163, n3000, n3003, n3004, Ng29161, n3005, Ng29160, n3006, Ng29159, n3008, n3007, n3009, Ng29158, n3010, Ng29157, n3011, Ng29156, n3013, n3016, n3017, Ng29153, n3018, Ng29152, n3019, Ng29151, n3021, n3020, n3022, Ng29150, n3023, Ng29149, n3024, Ng29148, n3026, n3029, n3030, Ng29145, n3031, Ng29144, n3032, Ng29143, n3034, n3033, n3035, Ng29142, n3036, Ng29141, n3037, Ng29140, n3039, n3042, n3043, Ng29137, n3044, Ng29136, n3045, Ng29135, n3047, n3046, n3048, Ng29134, n3049, Ng29133, n3050, Ng29132, n3051, Ng28308, n3052, Ng28307, n3053, Ng28306, n3055, n3056, Ng28305, n3057, Ng28304, n3058, Ng28303, n3060, n3061, Ng28302, n3062, Ng28301, n3063, Ng28300, n3064, Ng28299, n3065, Ng28298, n3066, Ng28297, n3067, Ng28296, n3068, Ng28295, n3069, Ng28294, n3071, n3072, Ng28293, n3073, Ng28292, n3074, Ng28291, n3076, n3077, Ng28290, n3078, Ng28289, n3079, Ng28288, n3080, Ng28287, n3081, Ng28286, n3082, Ng28285, n3083, Ng28282, n3084, Ng28281, n3085, Ng28280, n3087, n3088, Ng28279, n3089, Ng28278, n3090, Ng28277, n3092, n3093, Ng28276, n3094, Ng28275, n3095, Ng28274, n3096, Ng28273, n3097, Ng28272, n3098, Ng28271, n3099, Ng28270, n3100, Ng28269, n3101, Ng28268, n3103, n3104, Ng28267, n3105, Ng28266, n3106, Ng28265, n3108, n3109, Ng28264, n3110, Ng28263, n3111, Ng28262, n3112, Ng28261, n3113, Ng28260, n3114, Ng28259, n3115, Ng28256, n3116, Ng28255, n3117, Ng28254, n3119, n3120, Ng28253, n3121, Ng28252, n3122, Ng28251, n3124, n3125, Ng28250, n3126, Ng28249, n3127, Ng28248, n3128, Ng28247, n3129, Ng28246, n3130, Ng28245, n3131, Ng28244, n3132, Ng28243, n3133, Ng28242, n3135, n3136, Ng28241, n3137, Ng28240, n3138, Ng28239, n3140, n3141, Ng28238, n3142, Ng28237, n3143, Ng28236, n3144, Ng28235, n3145, Ng28234, n3146, Ng28233, n3147, Ng28230, n3148, Ng28229, n3149, Ng28228, n3151, n3152, Ng28227, n3153, Ng28226, n3154, Ng28225, n3156, n3157, Ng28224, n3158, Ng28223, n3159, Ng28222, n3160, Ng28221, n3161, Ng28220, n3162, Ng28219, n3163, Ng28218, n3164, Ng28217, n3165, Ng28216, n3167, n3168, Ng28215, n3169, Ng28214, n3170, Ng28213, n3172, n3173, Ng28212, n3174, Ng28211, n3175, Ng28210, n3176, Ng28209, n3177, Ng28208, n3178, Ng28207, n3179, Ng27713, n3180, Ng27712, n3181, Ng27711, n3182, Ng27710, n3183, Ng27709, n3184, Ng27708, n3185, Ng27705, n3186, Ng27704, n3187, Ng27703, n3188, Ng27702, n3189, Ng27701, n3190, Ng27700, n3191, Ng27697, n3192, Ng27696, n3193, Ng27695, n3194, Ng27694, n3195, Ng27693, n3196, Ng27692, n3197, Ng27689, n3198, Ng27688, n3199, Ng27687, n3200, Ng27686, n3201, Ng27685, n3202, Ng27684, n3203, Ng27235, n3204, Ng27234, n3205, Ng27233, n3206, Ng27232, n3207, Ng27231, n3208, Ng27230, n3209, Ng27226, n3210, Ng27225, n3211, Ng27224, n3212, Ng27223, n3213, Ng27222, n3214, Ng27221, n3215, Ng27211, n3216, Ng27210, n3217, Ng27209, n3218, Ng27208, n3219, Ng27207, n3220, Ng27206, n3221, Ng27196, n3222, Ng27195, n3223, Ng27194, n3224, Ng27193, n3225, Ng27192, n3226, Ng27191, n3227, Ng26753, n3228, Ng26752, n3229, Ng26751, n3230, Ng26748, n3231, Ng26745, n3232, Ng26744, n3233, Ng26743, n3234, Ng26741, n3235, Ng26740, n3236, Ng26739, n3237, Ng26738, n3238, Ng26737, n3239, Ng26736, n3240, Ng26735, n3241, Ng26734, n3242, Ng26733, n3243, Ng26732, n3244, Ng26731, n3245, Ng26730, n3246, Ng26728, n3247, Ng26727, n3248, Ng26726, n3249, Ng26724, n3250, Ng26723, n3251, Ng26722, n3252, Ng26721, n3253, Ng26720, n3254, Ng26719, n3255, Ng26718, n3256, Ng26717, n3257, Ng26716, n3258, Ng26715, n3259, Ng26714, n3260, Ng26713, n3261, Ng26711, n3262, Ng26710, n3263, Ng26709, n3264, Ng26707, n3265, Ng26706, n3266, Ng26705, n3267, Ng26704, n3268, Ng26703, n3269, Ng26702, n3270, Ng26701, n3271, Ng26700, n3272, Ng26699, n3273, Ng26698, n3274, Ng26697, n3275, Ng26696, n3276, Ng26694, n3277, Ng26693, n3278, Ng26692, n3279, Ng26690, n3280, Ng26689, n3281, Ng26688, n3282, Ng26687, n3283, Ng26686, n3284, Ng26685, n3285, Ng26684, n3286, Ng26683, n3287, Ng26682, n3288, Ng26681, n3289, Ng26680, n3290, Ng26679, n3291, Ng26017, n3292, Ng26016, n3293, Ng26015, n3294, Ng26014, n3295, Ng26013, n3296, Ng26012, n3297, Ng26011, n3298, Ng26010, n3299, Ng26008, n3300, Ng26007, n3301, Ng26006, n3302, Ng26005, n3303, Ng26004, n3304, Ng26003, n3305, Ng26002, n3306, Ng26001, n3307, Ng25999, n3308, Ng25998, n3309, Ng25997, n3310, Ng25996, n3311, Ng25995, n3312, Ng25994, n3313, Ng25993, n3314, Ng25992, n3315, Ng25990, n3316, Ng25989, n3317, Ng25988, n3318, Ng25987, n3319, Ng25986, n3320, Ng25985, n3321, Ng25984, n3322, Ng25983, n3323, n3324, Ng25172, n3325, Ng25171, n3326, Ng25170, n3327, Ng25169, n3328, Ng25168, n3329, Ng25167, n3330, Ng25166, n3331, Ng25165, n3332, Ng25164, n3333, Ng25161, n3334, Ng25160, n3335, Ng25159, n3336, Ng25158, n3337, Ng25157, n3338, Ng25156, n3339, Ng25155, n3340, Ng25154, n3341, Ng25153, n3342, Ng25150, n3343, Ng25149, n3344, Ng25148, n3345, Ng25147, n3346, Ng25146, n3347, Ng25145, n3348, Ng25144, n3349, Ng25143, n3350, Ng25142, n3351, Ng25139, n3352, Ng25138, n3353, Ng25137, n3354, Ng25136, n3355, Ng25135, n3356, Ng25134, n3357, Ng25133, n3358, Ng25132, n3359, Ng25131, n3360, Ng24417, n3361, Ng24416, n3362, Ng24415, n3363, Ng24414, n3364, Ng24413, n3365, Ng24412, n3366, Ng24411, n3367, Ng24410, n3368, Ng24409, n3369, Ng24408, n3370, Ng24407, n3371, Ng24406, n3372, Ng24405, n3373, Ng24404, n3374, Ng24403, n3375, Ng24402, n3376, Ng24401, n3377, Ng24400, n3378, Ng24399, n3379, Ng24398, n3380, Ng24397, n3381, Ng24396, n3382, Ng24395, n3383, Ng24394, n3384, Ng24393, n3385, Ng24392, n3386, Ng24391, n3387, Ng24390, n3388, Ng24389, n3389, Ng24388, n3390, Ng24387, n3391, Ng24386, n3392, Ng24385, n3393, Ng24384, n3394, Ng24383, n3395, Ng24382, n3396, Ng24376, n3397, Ng24375, n3398, Ng24374, n3399, Ng24373, n3400, Ng24372, n3401, Ng24371, n3402, Ng24370, n3403, Ng24369, n3404, Ng24368, n3405, Ng24367, n3406, Ng24366, n3407, Ng24365, n3408, Ng24364, n3409, Ng24363, n3410, Ng24362, n3411, Ng24361, n3412, Ng24360, n3413, Ng24359, n3414, Ng24358, n3415, Ng24357, n3416, Ng24356, n3417, Ng24355, n3418, Ng24354, n3419, Ng24353, n3420, Ng24352, n3421, Ng24351, n3422, Ng24350, n3423, Ng24349, n3424, Ng24348, n3425, Ng24347, n3426, Ng24346, n3427, Ng24345, n3428, Ng24344, n3429, Ng24343, n3430, Ng24342, n3431, Ng24341, n3432, Ng24335, n3433, Ng24334, n3434, Ng24333, n3435, Ng24332, n3436, Ng24331, n3437, Ng24330, n3438, Ng24329, n3439, Ng24328, n3440, Ng24327, n3441, Ng24326, n3442, Ng24325, n3443, Ng24324, n3444, Ng24323, n3445, Ng24322, n3446, Ng24321, n3447, Ng24320, n3448, Ng24319, n3449, Ng24318, n3450, Ng24317, n3451, Ng24316, n3452, Ng24315, n3453, Ng24314, n3454, Ng24313, n3455, Ng24312, n3456, Ng24311, n3457, Ng24310, n3458, Ng24309, n3459, Ng24308, n3460, Ng24307, n3461, Ng24306, n3462, Ng24305, n3463, Ng24304, n3464, Ng24303, n3465, Ng24302, n3466, Ng24301, n3467, Ng24300, n3468, Ng24294, n3469, Ng24293, n3470, Ng24292, n3471, Ng24291, n3472, Ng24290, n3473, Ng24289, n3474, Ng24288, n3475, Ng24287, n3476, Ng24286, n3477, Ng24285, n3478, Ng24284, n3479, Ng24283, n3480, Ng24282, n3481, Ng24281, n3482, Ng24280, n3483, Ng24279, n3484, Ng24278, n3485, Ng24277, n3486, Ng24276, n3487, Ng24275, n3488, Ng24274, n3489, Ng24273, n3490, Ng24272, n3491, Ng24271, n3492, Ng24270, n3493, Ng24269, n3494, Ng24268, n3495, Ng24267, n3496, Ng24266, n3497, Ng24265, n3498, Ng24264, n3499, Ng24263, n3500, Ng24262, n3501, Ng24261, n3502, Ng24260, n3503, Ng24259, n3504, Ng23316, n3505, Ng23314, n3506, Ng23313, n3507, Ng23312, n3508, Ng23311, n3509, Ng23310, n3510, Ng23309, n3511, Ng23308, n3512, Ng23307, n3513, Ng23306, n3514, Ng23305, n3515, Ng23304, n3516, Ng23303, n3517, Ng23302, n3518, Ng23301, n3519, Ng23300, n3520, Ng23299, n3521, Ng23298, n3522, Ng23297, n3523, Ng23296, n3524, Ng23295, n3525, Ng23294, n3526, Ng23293, n3527, Ng23292, n3528, Ng23291, n3529, Ng23290, n3530, Ng23289, n3531, Ng23288, n3532, Ng23287, n3533, Ng23286, n3534, Ng23285, n3535, Ng23284, n3536, Ng23283, n3537, Ng23282, n3538, Ng23281, n3539, Ng23280, n3540, Ng23279, n3541, Ng23278, n3542, Ng23277, n3543, Ng23276, n3544, Ng23273, n3545, Ng23272, n3546, Ng23271, n3547, Ng23270, n3548, Ng23269, n3549, Ng23268, n3550, Ng23267, n3551, Ng23266, n3552, Ng23265, n3553, Ng23264, n3554, Ng23263, n3555, Ng23262, n3556, Ng23261, n3557, Ng23260, n3558, Ng23259, n3559, Ng23258, n3560, Ng23257, n3561, Ng23256, n3562, Ng23255, n3563, Ng23254, n3564, Ng23253, n3565, Ng23252, n3566, Ng23251, n3567, Ng23250, n3568, Ng23249, n3569, Ng23248, n3570, Ng23247, n3571, Ng23246, n3572, Ng23245, n3573, Ng23244, n3574, Ng23243, n3575, Ng23242, n3576, Ng23241, n3577, Ng23240, n3578, Ng23239, n3579, Ng23238, n3580, Ng23235, n3581, Ng23234, n3582, Ng23233, n3583, Ng23232, n3584, Ng23231, n3585, Ng23230, n3586, Ng23229, n3587, Ng23228, n3588, Ng23227, n3589, Ng23226, n3590, Ng23225, n3591, Ng23224, n3592, Ng23223, n3593, Ng23222, n3594, Ng23221, n3595, Ng23220, n3596, Ng23219, n3597, Ng23218, n3598, Ng23217, n3599, Ng23216, n3600, Ng23215, n3601, Ng23214, n3602, Ng23213, n3603, Ng23212, n3604, Ng23211, n3605, Ng23210, n3606, Ng23209, n3607, Ng23208, n3608, Ng23207, n3609, Ng23206, n3610, Ng23205, n3611, Ng23204, n3612, Ng23203, n3613, Ng23202, n3614, Ng23201, n3615, Ng23200, n3616, Ng23197, n3617, Ng23196, n3618, Ng23195, n3619, Ng23194, n3620, Ng23193, n3621, Ng23192, n3622, Ng23191, n3623, Ng23190, n3624, Ng23189, n3625, Ng23188, n3626, Ng23187, n3627, Ng23186, n3628, Ng23185, n3629, Ng23184, n3630, Ng23183, n3631, Ng23182, n3632, Ng23181, n3633, Ng23180, n3634, Ng23179, n3635, Ng23178, n3636, Ng23177, n3637, Ng23176, n3638, Ng23175, n3639, Ng23174, n3640, Ng23173, n3641, Ng23172, n3642, Ng23171, n3643, Ng23170, n3644, Ng23169, n3645, Ng23168, n3646, Ng23167, n3647, Ng23166, n3648, Ng23165, n3649, Ng23164, n3650, Ng23163, n3651, Ng23162, n3652, Ng21963, n3653, Ng21962, n3654, Ng21961, n3655, Ng21960, n3656, Ng21959, n3657, Ng21958, n3658, Ng21957, n3659, Ng21956, n3660, Ng21955, n3661, Ng21954, n3662, Ng21953, n3663, Ng21952, n3664, Ng21950, n3665, Ng21949, n3666, Ng21948, n3667, Ng21947, n3668, Ng20632, n3669, Ng20631, n3670, Ng20630, n3671, Ng20629, n3672, Ng20628, n3673, Ng20627, n3674, Ng20626, n3675, Ng20625, n3676, Ng20624, n3677, Ng20623, n3678, Ng20622, n3679, Ng20621, n3680, Ng20620, n3681, Ng20619, n3682, Ng20618, n3683, Ng20617, n3684, Ng20616, n3685, Ng20615, n3686, Ng20614, n3687, Ng20613, n3688, Ng20612, n3689, Ng20611, n3690, Ng20610, n3691, Ng20609, n3692, Ng20608, n3693, Ng20607, n3694, Ng20606, n3695, Ng20605, n3696, Ng20603, n3697, Ng20602, n3698, Ng20601, n3699, Ng20600, n3700, Ng20599, n3701, Ng20598, n3702, Ng20597, n3703, Ng20596, n3704, Ng20595, n3705, Ng20593, n3706, Ng20592, n3707, Ng20591, n3708, Ng20590, n3709, Ng20589, n3710, Ng20587, n3711, Ng20586, n3712, Ng20585, n3713, Ng20584, n3714, Ng20583, n3715, Ng20582, n3716, Ng20581, n3717, Ng20580, n3718, Ng20579, n3719, Ng20578, n3720, Ng20577, n3721, Ng20576, n3722, Ng20575, n3723, Ng20574, n3724, Ng20573, n3725, Ng20572, n3726, Ng20570, n3727, Ng20569, n3728, Ng20568, n3729, Ng20566, n3730, Ng20565, n3731, Ng20564, n3732, Ng20562, n3733, Ng20561, n3734, Ng20560, n3735, Ng20558, n3736, Ng20557, n3737, Ng20556, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3746, n3748, n3749, n3750, n3751, n3752, n3754, n3755, n3756, n3758, n3760, n3762, n3763, n3764, n3765, n3766, n3768, n3769, n3770, n3772, n3774, n3776, n3779, n3781, n3783, n3785, n3787, n3789, n3792, n3794, n3796, n3798, n3800, n3802, n3805, n3807, n3809, n3811, n3813, n3815, n3818, n3820, n3822, n3824, n3826, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3838, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3849, n3848, n3850, n3852, n3851, n3853, n3855, n3854, n3856, n3858, n3857, n3859, n3860, n3861, n3862, n3863, n3864, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3884, n3886, n3889, n3892, n3895, n3897, n3898, n3900, n3904, n3905, n3907, n3909, n3910, n3912, n3913, n3916, n3925, n3926, n3928, n3929, n3932, n3941, n3942, n3944, n3945, n3948, n3957, n3958, n3960, n3961, n3964, n3973, n3978, n3983, n3988, n3993, n3994, n3996, n3995, n3997, n3998, n4000, n3999, n4001, n4002, n4004, n4003, n4005, n4006, n4008, n4007, n4010, Ng23154, n4011, Ng27212, n4013, n4016, n4020, n4022, n4025, n4028, n4031, n4032, n4034, n4037, n4041, n4045, n4049, n4054, n4055, n4057, n4059, n4060, n4062, n4066, n4069, n4071, n4072, n4074, n4078, n4081, n4083, n4084, n4086, n4090, n4093, n4095, n4096, n4098, n4102, n4105, n4108, n4107, n4110, n4109, n4112, n4111, n4114, n4113, n4118, n4116, n4120, n4123, n4122, n4125, n4128, n4127, n4130, n4133, n4132, n4135, n4136, n4137, n4138, n4139, n4140, n4142, n4144, n4147, n4150, n4158, n4163, n4165, n4167, n4170, n4181, n4187, n4189, n4191, n4194, n4197, n4205, n4210, n4212, n4214, n4217, n4228, n4234, n4236, n4238, n4241, n4244, n4252, n4257, n4259, n4261, n4264, n4275, n4281, n4283, n4285, n4288, n4291, n4299, n4304, n4306, n4308, n4311, n4322, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4339, n4341, n4344, n4347, n4349, n4352, n4354, n4357, n4359, n4362, n4370, n4373, n4375, n4385, n4404, n4423, n4442, n4445, n4446, n4447, n4449, n4450, n4451, n4452, n4453, n4454, n4456, n4455, n4503, n4506, n4644, n4869, Ng20567, n4870, n4871, n4872, n4873, n4878, n4893, n4894, n4895, n4896, n4897, n4898, n4900, n4904, n4905, n4906, n4907;

reg Pg8021, Ng2817, Ng2933, Ng13457, Ng2883, Ng2888, Ng2896, Ng2892, Ng2903, Ng2900, Ng2908, Ng2912, Ng2917, Ng2924, Ng2920, Ng2984, Ng2985, Ng2929, Ng2879, Ng2934, Ng2935, Ng2938, Ng2941, Ng2944, Ng2947, Ng2953, Ng2956, Ng2959, Ng2962, Ng2963, Ng2966, Ng2969, Ng2972, Ng2975, Ng2978, Ng2981, Ng2874, Ng1506, Ng1501, Ng1496, Ng1491, Ng1486, Ng1481, Ng1476, Ng1471, Ng13439, Pg8251, Ng813, Pg4090, Ng809, Pg4323, Ng805, Pg4590, Ng801, Pg6225, Ng797, Pg6442, Ng793, Pg6895, Ng789, Pg7334, Ng785, Pg7519, Ng13423, Pg8249, Ng125, Pg4088, Ng121, Pg4321, Ng117, Pg8023, Ng113, Pg8175, Ng109, Pg3993, Ng105, Pg4200, Ng101, Pg4450, Ng97, Pg8096, Ng13407, Ng2200, Ng2195, Ng2190, Ng2185, Ng2180, Ng2175, Ng2170, Ng2165, Ng13455, Ng3210, Ng3211, Ng3084, Ng3085, Ng3086, Ng3087, Ng3091, Ng3092, Ng3093, Ng3094, Ng3095, Ng3096, Ng3097, Ng3098, Ng3099, Ng3100, Ng3101, Ng3102, Ng3103, Ng3104, Ng3105, Ng3106, Ng3107, Ng3108, Ng3155, Ng3158, Ng3161, Ng3164, Ng3167, Ng3170, Ng3173, Ng3176, Ng3179, Ng3182, Ng3185, Ng3088, Ng3191, Ng3128, Ng3126, Ng3125, Ng3123, Ng3120, Ng3110, Ng3139, Ng3135, Ng3147, Ng185, Ng130, Ng131, Ng129, Ng133, Ng134, Ng132, Ng142, Ng143, Ng141, Ng145, Ng146, Ng144, Ng148, Ng149, Ng147, Ng151, Ng152, Ng150, Ng154, Ng155, Ng153, Ng157, Ng158, Ng156, Ng160, Ng161, Ng159, Ng163, Ng164, Ng162, Ng169, Ng170, Ng168, Ng172, Ng173, Ng171, Ng175, Ng176, Ng174, Ng178, Ng179, Ng177, Ng186, Ng189, Ng192, Ng231, Ng234, Ng237, Ng195, Ng198, Ng201, Ng240, Ng243, Ng246, Ng204, Ng207, Ng210, Ng249, Ng252, Ng255, Ng213, Ng216, Ng219, Ng258, Ng261, Ng264, Ng222, Ng225, Ng228, Ng267, Ng270, Ng273, Ng92, Ng88, Ng83, Ng79, Ng74, Ng70, Ng65, Ng61, Ng56, Ng52, Ng11497, Ng11498, Ng11499, Ng11500, Ng11501, Ng11502, Ng11503, Ng11504, Ng11505, Ng11506, Ng11507, Ng11508, Ng408, Ng411, Ng414, Ng417, Ng420, Ng423, Ng427, Ng428, Ng426, Ng429, Ng432, Ng435, Ng438, Ng441, Ng444, Ng448, Ng449, Ng447, Ng312, Ng313, Ng314, Ng315, Ng316, Ng317, Ng318, Ng319, Ng320, Ng322, Ng323, Ng321, Ng403, Ng404, Ng402, Ng450, Ng451, Ng452, Ng453, Ng454, Ng279, Ng280, Ng281, Ng282, Ng283, Ng284, Ng285, Ng286, Ng287, Ng288, Ng289, Ng290, Ng291, Ng299, Ng305, Ng298, Ng342, Ng349, Ng350, Ng351, Ng352, Ng353, Ng357, Ng364, Ng365, Ng366, Ng367, Ng368, Ng372, Ng379, Ng380, Ng381, Ng382, Ng383, Ng387, Ng394, Ng395, Ng396, Ng397, Ng324, Ng554, Ng557, Ng510, Ng513, Ng523, Ng524, Ng564, Ng569, Ng570, Ng571, Ng572, Ng573, Ng574, Ng565, Ng566, Ng567, Ng568, Ng489, Ng486, Ng487, Ng488, Ng11512, Ng11515, Ng11516, Ng477, Ng478, Ng479, Ng480, Ng484, Ng464, Ng11517, Ng11513, Ng11514, Ng528, Ng535, Ng542, Ng543, Ng544, Ng548, Ng549, Ng8284, Ng558, Ng559, Ng576, Ng577, Ng575, Ng579, Ng580, Ng578, Ng582, Ng583, Ng581, Ng585, Ng586, Ng584, Ng587, Ng590, Ng593, Ng596, Ng599, Ng602, Ng614, Ng617, Ng620, Ng605, Ng608, Ng611, Ng490, Ng493, Ng496, Ng506, Ng507, Pg16297, Ng525, Ng529, Ng530, Ng531, Ng532, Ng533, Ng534, Ng536, Ng537, Ng538, Ng541, Ng630, Ng659, Ng640, Ng633, Ng653, Ng646, Ng660, Ng672, Ng666, Ng679, Ng686, Ng692, Ng699, Ng700, Ng698, Ng702, Ng703, Ng701, Ng705, Ng706, Ng704, Ng708, Ng709, Ng707, Ng711, Ng712, Ng710, Ng714, Ng715, Ng713, Ng717, Ng718, Ng716, Ng720, Ng721, Ng719, Ng723, Ng724, Ng722, Ng726, Ng727, Ng725, Ng729, Ng730, Ng728, Ng732, Ng733, Ng731, Ng735, Ng736, Ng734, Ng738, Ng739, Ng737, wire1612, wire1594, Ng853, Ng818, Ng819, Ng817, Ng821, Ng822, Ng820, Ng830, Ng831, Ng829, Ng833, Ng834, Ng832, Ng836, Ng837, Ng835, Ng839, Ng840, Ng838, Ng842, Ng843, Ng841, Ng845, Ng846, Ng844, Ng848, Ng849, Ng847, Ng851, Ng852, Ng850, Ng857, Ng858, Ng856, Ng860, Ng861, Ng859, Ng863, Ng864, Ng862, Ng866, Ng867, Ng865, Ng873, Ng876, Ng879, Ng918, Ng921, Ng924, Ng882, Ng885, Ng888, Ng927, Ng930, Ng933, Ng891, Ng894, Ng897, Ng936, Ng939, Ng942, Ng900, Ng903, Ng906, Ng945, Ng948, Ng951, Ng909, Ng912, Ng915, Ng954, Ng957, Ng960, Ng780, Ng776, Ng771, Ng767, Ng762, Ng758, Ng753, Ng749, Ng744, Ng740, Ng11524, Ng11525, Ng11526, Ng11527, Ng11528, Ng11529, Ng11530, Ng11531, Ng11532, Ng11533, Ng11534, Ng11535, Ng1095, Ng1098, Ng1101, Ng1104, Ng1107, Ng1110, Ng1114, Ng1115, Ng1113, Ng1116, Ng1119, Ng1122, Ng1125, Ng1128, Ng1131, Ng1135, Ng1136, Ng1134, Ng999, Ng1000, Ng1001, Ng1002, Ng1003, Ng1004, Ng1005, Ng1006, Ng1007, Ng1009, Ng1010, Ng1008, Ng1090, Ng1091, Ng1089, Ng1137, Ng1138, Ng1139, Ng1140, Ng1141, Ng966, Ng967, Ng968, Ng969, Ng970, Ng971, Ng972, Ng973, Ng974, Ng975, Ng976, Ng977, Ng978, Ng986, Ng992, Ng985, Ng1029, Ng1036, Ng1037, Ng1038, Ng1039, Ng1040, Ng1044, Ng1051, Ng1052, Ng1053, Ng1054, Ng1055, Ng1059, Ng1066, Ng1067, Ng1068, Ng1069, Ng1070, Ng1074, Ng1081, Ng1082, Ng1083, Ng1084, Ng1011, Ng1240, Ng1243, Ng1196, Ng1199, Ng1209, Ng1210, Ng1250, Ng1255, Ng1256, Ng1257, Ng1258, Ng1259, Ng1260, Ng1251, Ng1252, Ng1253, Ng1254, Ng1176, Ng1173, Ng1174, Ng1175, Ng11539, Ng11542, Ng11543, Ng1164, Ng1165, Ng1166, Ng1167, Ng1171, Ng1151, Ng11544, Ng11540, Ng11541, Ng1214, Ng1221, Ng1228, Ng1229, Ng1230, Ng1234, Ng1235, Ng8293, Ng1244, Ng1245, Ng1262, Ng1263, Ng1261, Ng1265, Ng1266, Ng1264, Ng1268, Ng1269, Ng1267, Ng1271, Ng1272, Ng1270, Ng1273, Ng1276, Ng1279, Ng1282, Ng1285, Ng1288, Ng1300, Ng1303, Ng1306, Ng1291, Ng1294, Ng1297, Ng1177, Ng1180, Ng1183, Ng1192, Ng1193, Pg16355, Ng1211, Ng1215, Ng1216, Ng1217, Ng1218, Ng1219, Ng1220, Ng1222, Ng1223, Ng1224, Ng1227, wire1605, wire1603, Ng1315, Ng1316, Ng1345, Ng1326, Ng1319, Ng1339, Ng1332, Ng1346, Ng1358, Ng1352, Ng1365, Ng1372, Ng1378, Ng1385, Ng1386, Ng1384, Ng1388, Ng1389, Ng1387, Ng1391, Ng1392, Ng1390, Ng1394, Ng1395, Ng1393, Ng1397, Ng1398, Ng1396, Ng1400, Ng1401, Ng1399, Ng1403, Ng1404, Ng1402, Ng1406, Ng1407, Ng1405, Ng1409, Ng1410, Ng1408, Ng1412, Ng1413, Ng1411, Ng1415, Ng1416, Ng1414, Ng1418, Ng1419, Ng1417, Ng1421, Ng1422, Ng1420, Ng1424, Ng1425, Ng1423, Ng1512, Ng1513, Ng1511, Ng1515, Ng1516, Ng1514, Ng1524, Ng1525, Ng1523, Ng1527, Ng1528, Ng1526, Ng1530, Ng1531, Ng1529, Ng1533, Ng1534, Ng1532, Ng1536, Ng1537, Ng1535, Ng1539, Ng1540, Ng1538, Ng1542, Ng1543, Ng1541, Ng1545, Ng1546, Ng1544, Ng1551, Ng1552, Ng1550, Ng1554, Ng1555, Ng1553, Ng1557, Ng1558, Ng1556, Ng1560, Ng1561, Ng1559, Ng1567, Ng1570, Ng1573, Ng1612, Ng1615, Ng1618, Ng1576, Ng1579, Ng1582, Ng1621, Ng1624, Ng1627, Ng1585, Ng1588, Ng1591, Ng1630, Ng1633, Ng1636, Ng1594, Ng1597, Ng1600, Ng1639, Ng1642, Ng1645, Ng1603, Ng1606, Ng1609, Ng1648, Ng1651, Ng1654, Ng1466, Ng1462, Ng1457, Ng1453, Ng1448, Ng1444, Ng1439, Ng1435, Ng1430, Ng1426, Ng11551, Ng11552, Ng11553, Ng11554, Ng11555, Ng11556, Ng11557, Ng11558, Ng11559, Ng11560, Ng11561, Ng11562, Ng1789, Ng1792, Ng1795, Ng1798, Ng1801, Ng1804, Ng1808, Ng1809, Ng1807, Ng1810, Ng1813, Ng1816, Ng1819, Ng1822, Ng1825, Ng1829, Ng1830, Ng1828, Ng1693, Ng1694, Ng1695, Ng1696, Ng1697, Ng1698, Ng1699, Ng1700, Ng1701, Ng1703, Ng1704, Ng1702, Ng1784, Ng1785, Ng1783, Ng1831, Ng1832, Ng1833, Ng1834, Ng1835, Ng1660, Ng1661, Ng1662, Ng1663, Ng1664, Ng1665, Ng1666, Ng1667, Ng1668, Ng1669, Ng1670, Ng1671, Ng1672, Ng1680, Ng1686, Ng1679, Ng1723, Ng1730, Ng1731, Ng1732, Ng1733, Ng1734, Ng1738, Ng1745, Ng1746, Ng1747, Ng1748, Ng1749, Ng1753, Ng1760, Ng1761, Ng1762, Ng1763, Ng1764, Ng1768, Ng1775, Ng1776, Ng1777, Ng1778, Ng1705, Ng1934, Ng1937, Ng1890, Ng1893, Ng1903, Ng1904, Ng1944, Ng1949, Ng1950, Ng1951, Ng1952, Ng1953, Ng1954, Ng1945, Ng1946, Ng1947, Ng1948, Ng1870, Ng1867, Ng1868, Ng1869, Ng11566, Ng11569, Ng11570, Ng1858, Ng1859, Ng1860, Ng1861, Ng1865, Ng1845, Ng11571, Ng11567, Ng11568, Ng1908, Ng1915, Ng1922, Ng1923, Ng1924, Ng1928, Ng1929, Ng8302, Ng1938, Ng1939, Ng1956, Ng1957, Ng1955, Ng1959, Ng1960, Ng1958, Ng1962, Ng1963, Ng1961, Ng1965, Ng1966, Ng1964, Ng1967, Ng1970, Ng1973, Ng1976, Ng1979, Ng1982, Ng1994, Ng1997, Ng2000, Ng1985, Ng1988, Ng1991, Ng1871, Ng1874, Ng1877, Ng1886, Ng1887, Pg16399, Ng1905, Ng1909, Ng1910, Ng1911, Ng1912, Ng1913, Ng1914, Ng1916, Ng1917, Ng1918, Ng1921, Ng2010, Ng2039, Ng2020, Ng2013, Ng2033, Ng2026, Ng2040, Ng2052, Ng2046, Ng2059, Ng2066, Ng2072, Ng2079, Ng2080, Ng2078, Ng2082, Ng2083, Ng2081, Ng2085, Ng2086, Ng2084, Ng2088, Ng2089, Ng2087, Ng2091, Ng2092, Ng2090, Ng2094, Ng2095, Ng2093, Ng2097, Ng2098, Ng2096, Ng2100, Ng2101, Ng2099, Ng2103, Ng2104, Ng2102, Ng2106, Ng2107, Ng2105, Ng2109, Ng2110, Ng2108, Ng2112, Ng2113, Ng2111, Ng2115, Ng2116, Ng2114, Ng2118, Ng2119, Ng2117, Ng2206, Ng2207, Ng2205, Ng2209, Ng2210, Ng2208, Ng2218, Ng2219, Ng2217, Ng2221, Ng2222, Ng2220, Ng2224, Ng2225, Ng2223, Ng2227, Ng2228, Ng2226, Ng2230, Ng2231, Ng2229, Ng2233, Ng2234, Ng2232, Ng2236, Ng2237, Ng2235, Ng2239, Ng2240, Ng2238, Ng2245, Ng2246, Ng2244, Ng2248, Ng2249, Ng2247, Ng2251, Ng2252, Ng2250, Ng2254, Ng2255, Ng2253, Ng2261, Ng2264, Ng2267, Ng2306, Ng2309, Ng2312, Ng2270, Ng2273, Ng2276, Ng2315, Ng2318, Ng2321, Ng2279, Ng2282, Ng2285, Ng2324, Ng2327, Ng2330, Ng2288, Ng2291, Ng2294, Ng2333, Ng2336, Ng2339, Ng2297, Ng2300, Ng2303, Ng2342, Ng2345, Ng2348, Ng2160, Ng2156, Ng2151, Ng2147, Ng2142, Ng2138, Ng2133, Ng2129, Ng2124, Ng2120, Ng2256, wire1609, Ng2257, Ng11578, Ng11579, Ng11580, Ng11581, Ng11582, Ng11583, Ng11584, Ng11585, Ng11586, Ng11587, Ng11588, Ng11589, Ng2483, Ng2486, Ng2489, Ng2492, Ng2495, Ng2498, Ng2502, Ng2503, Ng2501, Ng2504, Ng2507, Ng2510, Ng2513, Ng2516, Ng2519, Ng2523, Ng2524, Ng2522, Ng2387, Ng2388, Ng2389, Ng2390, Ng2391, Ng2392, Ng2393, Ng2394, Ng2395, Ng2397, Ng2398, Ng2396, Ng2478, Ng2479, Ng2477, Ng2525, Ng2526, Ng2527, Ng2528, Ng2529, Ng2354, Ng2355, Ng2356, Ng2357, Ng2358, Ng2359, Ng2360, Ng2361, Ng2362, Ng2363, Ng2364, Ng2365, Ng2366, Ng2374, Ng2380, Ng2373, Ng2417, Ng2424, Ng2425, Ng2426, Ng2427, Ng2428, Ng2432, Ng2439, Ng2440, Ng2441, Ng2442, Ng2443, Ng2447, Ng2454, Ng2455, Ng2456, Ng2457, Ng2458, Ng2462, Ng2469, Ng2470, Ng2471, Ng2472, Ng2399, Ng2628, Ng2631, Ng2584, Ng2587, Ng2597, Ng2598, Ng2638, Ng2643, Ng2644, Ng2645, Ng2646, Ng2647, Ng2648, Ng2639, Ng2640, Ng2641, Ng2642, Ng2564, Ng2561, Ng2562, Ng2563, Ng11593, Ng11596, Ng11597, Ng2552, Ng2553, Ng2554, Ng2555, Ng2559, Ng2539, Ng11598, Ng11594, Ng11595, Ng2602, Ng2609, Ng2616, Ng2617, Ng2618, Ng2622, Ng2623, Ng8311, Ng2632, Ng2633, Ng2650, Ng2651, Ng2649, Ng2653, Ng2654, Ng2652, Ng2656, Ng2657, Ng2655, Ng2659, Ng2660, Ng2658, Ng2661, Ng2664, Ng2667, Ng2670, Ng2673, Ng2676, Ng2688, Ng2691, Ng2694, Ng2679, Ng2682, Ng2685, Ng2565, Ng2568, Ng2571, Ng2580, Ng2581, Pg16437, Ng2599, Ng2603, Ng2604, Ng2605, Ng2606, Ng2607, Ng2608, Ng2610, Ng2611, Ng2612, Ng2615, Ng2704, Ng2733, Ng2714, Ng2707, Ng2727, Ng2720, Ng2734, Ng2746, Ng2740, Ng2753, Ng2760, Ng2766, Ng2773, Ng2774, Ng2772, Ng2776, Ng2777, Ng2775, Ng2779, Ng2780, Ng2778, Ng2782, Ng2783, Ng2781, Ng2785, Ng2786, Ng2784, Ng2788, Ng2789, Ng2787, Ng2791, Ng2792, Ng2790, Ng2794, Ng2795, Ng2793, Ng2797, Ng2798, Ng2796, Ng2800, Ng2801, Ng2799, Ng2803, Ng2804, Ng2802, Ng2806, Ng2807, Ng2805, Ng2809, Ng2810, Ng2808, Ng2812, Ng2813, Ng2811, Ng3054, Ng3079, Ng13475, Ng3043, Ng3044, Ng3045, Ng3046, Ng3047, Ng3048, Ng3049, Ng3050, Ng3051, Ng3052, Ng3053, Ng3055, Ng3056, Ng3057, Ng3058, Ng3059, Ng3060, Ng3061, Ng3062, Ng3063, Ng3064, Ng3065, Ng3066, Ng3067, Ng3068, Ng3069, Ng3070, Ng3071, Ng3072, Ng3073, Ng3074, Ng3075, Ng3076, Ng3077, Ng3078, Ng2997, Ng2993, Ng2998, Ng3006, Ng3002, Ng3013, Ng3010, Ng3024, Ng3018, Ng3028, Ng3036, Ng3032, Pg5388, Ng2986, Ng2987, Pg8275, Pg8274, Pg8273, Pg8272, Pg8268, Pg8269, Pg8270, Pg8271, Ng3083, Pg8267, Ng2992, Pg8266, Pg8265, Pg8264, Pg8262, Pg8263, Pg8260, Pg8261, Pg8259, Ng2990, Ng2991, Pg8258;

always  @(posedge PCLK)
	Pg8021<=Pg51;

 always  @(posedge PCLK)
	Ng2817<=Ng20571;

 always  @(posedge PCLK)
	Ng2933<=Ng20588;

 always  @(posedge PCLK)
	Ng13457<=Ng21951;

 always  @(posedge PCLK)
	Ng2883<=Ng23315;

 always  @(posedge PCLK)
	Ng2888<=Ng24423;

 always  @(posedge PCLK)
	Ng2896<=Ng25175;

 always  @(posedge PCLK)
	Ng2892<=Ng26019;

 always  @(posedge PCLK)
	Ng2903<=Ng26747;

 always  @(posedge PCLK)
	Ng2900<=Ng27237;

 always  @(posedge PCLK)
	Ng2908<=Ng27715;

 always  @(posedge PCLK)
	Ng2912<=Ng24424;

 always  @(posedge PCLK)
	Ng2917<=Ng25174;

 always  @(posedge PCLK)
	Ng2924<=Ng26020;

 always  @(posedge PCLK)
	Ng2920<=Ng26746;

 always  @(posedge PCLK)
	Ng2984<=Ng19061;

 always  @(posedge PCLK)
	Ng2985<=Ng19060;

 always  @(posedge PCLK)
	Ng2929<=Pg8021;

 always  @(posedge PCLK)
	Ng2879<=Ng16494;

 always  @(posedge PCLK)
	Ng2934<=Pg3212;

 always  @(posedge PCLK)
	Ng2935<=Pg3228;

 always  @(posedge PCLK)
	Ng2938<=Pg3227;

 always  @(posedge PCLK)
	Ng2941<=Pg3226;

 always  @(posedge PCLK)
	Ng2944<=Pg3225;

 always  @(posedge PCLK)
	Ng2947<=Pg3224;

 always  @(posedge PCLK)
	Ng2953<=Pg3223;

 always  @(posedge PCLK)
	Ng2956<=Pg3222;

 always  @(posedge PCLK)
	Ng2959<=Pg3221;

 always  @(posedge PCLK)
	Ng2962<=Pg3232;

 always  @(posedge PCLK)
	Ng2963<=Pg3220;

 always  @(posedge PCLK)
	Ng2966<=Pg3219;

 always  @(posedge PCLK)
	Ng2969<=Pg3218;

 always  @(posedge PCLK)
	Ng2972<=Pg3217;

 always  @(posedge PCLK)
	Ng2975<=Pg3216;

 always  @(posedge PCLK)
	Ng2978<=Pg3215;

 always  @(posedge PCLK)
	Ng2981<=Pg3214;

 always  @(posedge PCLK)
	Ng2874<=Pg3213;

 always  @(posedge PCLK)
	Ng1506<=Ng20572;

 always  @(posedge PCLK)
	Ng1501<=Ng20573;

 always  @(posedge PCLK)
	Ng1496<=Ng20574;

 always  @(posedge PCLK)
	Ng1491<=Ng20575;

 always  @(posedge PCLK)
	Ng1486<=Ng20576;

 always  @(posedge PCLK)
	Ng1481<=Ng20577;

 always  @(posedge PCLK)
	Ng1476<=Ng20578;

 always  @(posedge PCLK)
	Ng1471<=Ng20579;

 always  @(posedge PCLK)
	Ng13439<=Ng23313;

 always  @(posedge PCLK)
	Pg8251<=Ng21960;

 always  @(posedge PCLK)
	Ng813<=Pg8251;

 always  @(posedge PCLK)
	Pg4090<=Ng21961;

 always  @(posedge PCLK)
	Ng809<=Pg4090;

 always  @(posedge PCLK)
	Pg4323<=Ng21962;

 always  @(posedge PCLK)
	Ng805<=Pg4323;

 always  @(posedge PCLK)
	Pg4590<=Ng21963;

 always  @(posedge PCLK)
	Ng801<=Pg4590;

 always  @(posedge PCLK)
	Pg6225<=Ng21947;

 always  @(posedge PCLK)
	Ng797<=Pg6225;

 always  @(posedge PCLK)
	Pg6442<=Ng21948;

 always  @(posedge PCLK)
	Ng793<=Pg6442;

 always  @(posedge PCLK)
	Pg6895<=Ng21949;

 always  @(posedge PCLK)
	Ng789<=Pg6895;

 always  @(posedge PCLK)
	Pg7334<=Ng21950;

 always  @(posedge PCLK)
	Ng785<=Pg7334;

 always  @(posedge PCLK)
	Pg7519<=Ng23312;

 always  @(posedge PCLK)
	Ng13423<=Pg7519;

 always  @(posedge PCLK)
	Pg8249<=Ng21952;

 always  @(posedge PCLK)
	Ng125<=Pg8249;

 always  @(posedge PCLK)
	Pg4088<=Ng21953;

 always  @(posedge PCLK)
	Ng121<=Pg4088;

 always  @(posedge PCLK)
	Pg4321<=Ng21954;

 always  @(posedge PCLK)
	Ng117<=Pg4321;

 always  @(posedge PCLK)
	Pg8023<=Ng21955;

 always  @(posedge PCLK)
	Ng113<=Pg8023;

 always  @(posedge PCLK)
	Pg8175<=Ng21956;

 always  @(posedge PCLK)
	Ng109<=Pg8175;

 always  @(posedge PCLK)
	Pg3993<=Ng21957;

 always  @(posedge PCLK)
	Ng105<=Pg3993;

 always  @(posedge PCLK)
	Pg4200<=Ng21958;

 always  @(posedge PCLK)
	Ng101<=Pg4200;

 always  @(posedge PCLK)
	Pg4450<=Ng21959;

 always  @(posedge PCLK)
	Ng97<=Pg4450;

 always  @(posedge PCLK)
	Pg8096<=Ng23316;

 always  @(posedge PCLK)
	Ng13407<=Pg8096;

 always  @(posedge PCLK)
	Ng2200<=Ng20587;

 always  @(posedge PCLK)
	Ng2195<=Ng20585;

 always  @(posedge PCLK)
	Ng2190<=Ng20586;

 always  @(posedge PCLK)
	Ng2185<=Ng20584;

 always  @(posedge PCLK)
	Ng2180<=Ng20583;

 always  @(posedge PCLK)
	Ng2175<=Ng20582;

 always  @(posedge PCLK)
	Ng2170<=Ng20581;

 always  @(posedge PCLK)
	Ng2165<=Ng20580;

 always  @(posedge PCLK)
	Ng13455<=Ng23314;

 always  @(posedge PCLK)
	Ng3210<=Ng20630;

 always  @(posedge PCLK)
	Ng3211<=Ng20631;

 always  @(posedge PCLK)
	Ng3084<=Ng20632;

 always  @(posedge PCLK)
	Ng3085<=Ng20609;

 always  @(posedge PCLK)
	Ng3086<=Ng20610;

 always  @(posedge PCLK)
	Ng3087<=Ng20611;

 always  @(posedge PCLK)
	Ng3091<=Ng20612;

 always  @(posedge PCLK)
	Ng3092<=Ng20613;

 always  @(posedge PCLK)
	Ng3093<=Ng20614;

 always  @(posedge PCLK)
	Ng3094<=Ng20615;

 always  @(posedge PCLK)
	Ng3095<=Ng20616;

 always  @(posedge PCLK)
	Ng3096<=Ng20617;

 always  @(posedge PCLK)
	Ng3097<=Ng26751;

 always  @(posedge PCLK)
	Ng3098<=Ng26752;

 always  @(posedge PCLK)
	Ng3099<=Ng26753;

 always  @(posedge PCLK)
	Ng3100<=Ng29163;

 always  @(posedge PCLK)
	Ng3101<=Ng29164;

 always  @(posedge PCLK)
	Ng3102<=Ng29165;

 always  @(posedge PCLK)
	Ng3103<=Ng30120;

 always  @(posedge PCLK)
	Ng3104<=Ng30121;

 always  @(posedge PCLK)
	Ng3105<=Ng30122;

 always  @(posedge PCLK)
	Ng3106<=Ng30941;

 always  @(posedge PCLK)
	Ng3107<=Ng30942;

 always  @(posedge PCLK)
	Ng3108<=Ng30943;

 always  @(posedge PCLK)
	Ng3155<=Ng20618;

 always  @(posedge PCLK)
	Ng3158<=Ng20619;

 always  @(posedge PCLK)
	Ng3161<=Ng20620;

 always  @(posedge PCLK)
	Ng3164<=Ng20621;

 always  @(posedge PCLK)
	Ng3167<=Ng20622;

 always  @(posedge PCLK)
	Ng3170<=Ng20623;

 always  @(posedge PCLK)
	Ng3173<=Ng20624;

 always  @(posedge PCLK)
	Ng3176<=Ng20625;

 always  @(posedge PCLK)
	Ng3179<=Ng20626;

 always  @(posedge PCLK)
	Ng3182<=Ng20627;

 always  @(posedge PCLK)
	Ng3185<=Ng20628;

 always  @(posedge PCLK)
	Ng3088<=Ng20629;

 always  @(posedge PCLK)
	Ng3191<=Pg24734;

 always  @(posedge PCLK)
	Ng3128<=Ng29166;

 always  @(posedge PCLK)
	Ng3126<=wire1521;

 always  @(posedge PCLK)
	Ng3125<=Ng28696;

 always  @(posedge PCLK)
	Ng3123<=Ng28313;

 always  @(posedge PCLK)
	Ng3120<=Pg26104;

 always  @(posedge PCLK)
	Ng3110<=Pg25435;

 always  @(posedge PCLK)
	Ng3139<=Pg27380;

 always  @(posedge PCLK)
	Ng3135<=Pg26149;

 always  @(posedge PCLK)
	Ng3147<=Pg26135;

 always  @(posedge PCLK)
	Ng185<=Ng29656;

 always  @(posedge PCLK)
	Ng130<=Ng24259;

 always  @(posedge PCLK)
	Ng131<=Ng24260;

 always  @(posedge PCLK)
	Ng129<=Ng24261;

 always  @(posedge PCLK)
	Ng133<=Ng24262;

 always  @(posedge PCLK)
	Ng134<=Ng24263;

 always  @(posedge PCLK)
	Ng132<=Ng24264;

 always  @(posedge PCLK)
	Ng142<=Ng24265;

 always  @(posedge PCLK)
	Ng143<=Ng24266;

 always  @(posedge PCLK)
	Ng141<=Ng24267;

 always  @(posedge PCLK)
	Ng145<=Ng24268;

 always  @(posedge PCLK)
	Ng146<=Ng24269;

 always  @(posedge PCLK)
	Ng144<=Ng24270;

 always  @(posedge PCLK)
	Ng148<=Ng24271;

 always  @(posedge PCLK)
	Ng149<=Ng24272;

 always  @(posedge PCLK)
	Ng147<=Ng24273;

 always  @(posedge PCLK)
	Ng151<=Ng24274;

 always  @(posedge PCLK)
	Ng152<=Ng24275;

 always  @(posedge PCLK)
	Ng150<=Ng24276;

 always  @(posedge PCLK)
	Ng154<=Ng24277;

 always  @(posedge PCLK)
	Ng155<=Ng24278;

 always  @(posedge PCLK)
	Ng153<=Ng24279;

 always  @(posedge PCLK)
	Ng157<=Ng24280;

 always  @(posedge PCLK)
	Ng158<=Ng24281;

 always  @(posedge PCLK)
	Ng156<=Ng24282;

 always  @(posedge PCLK)
	Ng160<=Ng24283;

 always  @(posedge PCLK)
	Ng161<=Ng24284;

 always  @(posedge PCLK)
	Ng159<=Ng24285;

 always  @(posedge PCLK)
	Ng163<=Ng24286;

 always  @(posedge PCLK)
	Ng164<=Ng24287;

 always  @(posedge PCLK)
	Ng162<=Ng24288;

 always  @(posedge PCLK)
	Ng169<=Ng26679;

 always  @(posedge PCLK)
	Ng170<=Ng26680;

 always  @(posedge PCLK)
	Ng168<=Ng26681;

 always  @(posedge PCLK)
	Ng172<=Ng26682;

 always  @(posedge PCLK)
	Ng173<=Ng26683;

 always  @(posedge PCLK)
	Ng171<=Ng26684;

 always  @(posedge PCLK)
	Ng175<=Ng26685;

 always  @(posedge PCLK)
	Ng176<=Ng26686;

 always  @(posedge PCLK)
	Ng174<=Ng26687;

 always  @(posedge PCLK)
	Ng178<=Ng26688;

 always  @(posedge PCLK)
	Ng179<=Ng26689;

 always  @(posedge PCLK)
	Ng177<=Ng26690;

 always  @(posedge PCLK)
	Ng186<=Ng30506;

 always  @(posedge PCLK)
	Ng189<=Ng30507;

 always  @(posedge PCLK)
	Ng192<=Ng30508;

 always  @(posedge PCLK)
	Ng231<=Ng30842;

 always  @(posedge PCLK)
	Ng234<=Ng30843;

 always  @(posedge PCLK)
	Ng237<=Ng30844;

 always  @(posedge PCLK)
	Ng195<=Ng30836;

 always  @(posedge PCLK)
	Ng198<=Ng30837;

 always  @(posedge PCLK)
	Ng201<=Ng30838;

 always  @(posedge PCLK)
	Ng240<=Ng30845;

 always  @(posedge PCLK)
	Ng243<=Ng30846;

 always  @(posedge PCLK)
	Ng246<=Ng30847;

 always  @(posedge PCLK)
	Ng204<=Ng30509;

 always  @(posedge PCLK)
	Ng207<=Ng30510;

 always  @(posedge PCLK)
	Ng210<=Ng30511;

 always  @(posedge PCLK)
	Ng249<=Ng30515;

 always  @(posedge PCLK)
	Ng252<=Ng30516;

 always  @(posedge PCLK)
	Ng255<=Ng30517;

 always  @(posedge PCLK)
	Ng213<=Ng30512;

 always  @(posedge PCLK)
	Ng216<=Ng30513;

 always  @(posedge PCLK)
	Ng219<=Ng30514;

 always  @(posedge PCLK)
	Ng258<=Ng30518;

 always  @(posedge PCLK)
	Ng261<=Ng30519;

 always  @(posedge PCLK)
	Ng264<=Ng30520;

 always  @(posedge PCLK)
	Ng222<=Ng30839;

 always  @(posedge PCLK)
	Ng225<=Ng30840;

 always  @(posedge PCLK)
	Ng228<=Ng30841;

 always  @(posedge PCLK)
	Ng267<=Ng30848;

 always  @(posedge PCLK)
	Ng270<=Ng30849;

 always  @(posedge PCLK)
	Ng273<=Ng30850;

 always  @(posedge PCLK)
	Ng92<=Ng25983;

 always  @(posedge PCLK)
	Ng88<=Ng26678;

 always  @(posedge PCLK)
	Ng83<=Ng27189;

 always  @(posedge PCLK)
	Ng79<=Ng27683;

 always  @(posedge PCLK)
	Ng74<=Ng28206;

 always  @(posedge PCLK)
	Ng70<=Ng28673;

 always  @(posedge PCLK)
	Ng65<=Ng29131;

 always  @(posedge PCLK)
	Ng61<=Ng29413;

 always  @(posedge PCLK)
	Ng56<=Ng29627;

 always  @(posedge PCLK)
	Ng52<=Ng29794;

 always  @(posedge PCLK)
	Ng11497<=Ng28207;

 always  @(posedge PCLK)
	Ng11498<=Ng28208;

 always  @(posedge PCLK)
	Ng11499<=Ng28209;

 always  @(posedge PCLK)
	Ng11500<=Ng28210;

 always  @(posedge PCLK)
	Ng11501<=Ng28211;

 always  @(posedge PCLK)
	Ng11502<=Ng28212;

 always  @(posedge PCLK)
	Ng11503<=Ng28213;

 always  @(posedge PCLK)
	Ng11504<=Ng28214;

 always  @(posedge PCLK)
	Ng11505<=Ng28215;

 always  @(posedge PCLK)
	Ng11506<=Ng28216;

 always  @(posedge PCLK)
	Ng11507<=Ng28217;

 always  @(posedge PCLK)
	Ng11508<=Ng28218;

 always  @(posedge PCLK)
	Ng408<=Ng29414;

 always  @(posedge PCLK)
	Ng411<=Ng29415;

 always  @(posedge PCLK)
	Ng414<=Ng29416;

 always  @(posedge PCLK)
	Ng417<=Ng29631;

 always  @(posedge PCLK)
	Ng420<=Ng29632;

 always  @(posedge PCLK)
	Ng423<=Ng29633;

 always  @(posedge PCLK)
	Ng427<=Ng29417;

 always  @(posedge PCLK)
	Ng428<=Ng29418;

 always  @(posedge PCLK)
	Ng426<=Ng29419;

 always  @(posedge PCLK)
	Ng429<=Ng27684;

 always  @(posedge PCLK)
	Ng432<=Ng27685;

 always  @(posedge PCLK)
	Ng435<=Ng27686;

 always  @(posedge PCLK)
	Ng438<=Ng27687;

 always  @(posedge PCLK)
	Ng441<=Ng27688;

 always  @(posedge PCLK)
	Ng444<=Ng27689;

 always  @(posedge PCLK)
	Ng448<=Ng28674;

 always  @(posedge PCLK)
	Ng449<=Ng28675;

 always  @(posedge PCLK)
	Ng447<=Ng28676;

 always  @(posedge PCLK)
	Ng312<=Ng29795;

 always  @(posedge PCLK)
	Ng313<=Ng29796;

 always  @(posedge PCLK)
	Ng314<=Ng29797;

 always  @(posedge PCLK)
	Ng315<=Ng30851;

 always  @(posedge PCLK)
	Ng316<=Ng30852;

 always  @(posedge PCLK)
	Ng317<=Ng30853;

 always  @(posedge PCLK)
	Ng318<=Ng30710;

 always  @(posedge PCLK)
	Ng319<=Ng30711;

 always  @(posedge PCLK)
	Ng320<=Ng30712;

 always  @(posedge PCLK)
	Ng322<=Ng29628;

 always  @(posedge PCLK)
	Ng323<=Ng29629;

 always  @(posedge PCLK)
	Ng321<=Ng29630;

 always  @(posedge PCLK)
	Ng403<=Ng27191;

 always  @(posedge PCLK)
	Ng404<=Ng27192;

 always  @(posedge PCLK)
	Ng402<=Ng27193;

 always  @(posedge PCLK)
	Ng450<=Ng11509;

 always  @(posedge PCLK)
	Ng451<=Ng450;

 always  @(posedge PCLK)
	Ng452<=Ng11510;

 always  @(posedge PCLK)
	Ng453<=Ng452;

 always  @(posedge PCLK)
	Ng454<=Ng11511;

 always  @(posedge PCLK)
	Ng279<=Ng454;

 always  @(posedge PCLK)
	Ng280<=Ng11491;

 always  @(posedge PCLK)
	Ng281<=Ng280;

 always  @(posedge PCLK)
	Ng282<=Ng11492;

 always  @(posedge PCLK)
	Ng283<=Ng282;

 always  @(posedge PCLK)
	Ng284<=Ng11493;

 always  @(posedge PCLK)
	Ng285<=Ng284;

 always  @(posedge PCLK)
	Ng286<=Ng11494;

 always  @(posedge PCLK)
	Ng287<=Ng286;

 always  @(posedge PCLK)
	Ng288<=Ng11495;

 always  @(posedge PCLK)
	Ng289<=Ng288;

 always  @(posedge PCLK)
	Ng290<=Ng13407;

 always  @(posedge PCLK)
	Ng291<=Ng290;

 always  @(posedge PCLK)
	Ng299<=Ng19012;

 always  @(posedge PCLK)
	Ng305<=Ng23148;

 always  @(posedge PCLK)
	Ng298<=Ng27190;

 always  @(posedge PCLK)
	Ng342<=Ng11497;

 always  @(posedge PCLK)
	Ng349<=Ng342;

 always  @(posedge PCLK)
	Ng350<=Ng11498;

 always  @(posedge PCLK)
	Ng351<=Ng350;

 always  @(posedge PCLK)
	Ng352<=Ng11499;

 always  @(posedge PCLK)
	Ng353<=Ng352;

 always  @(posedge PCLK)
	Ng357<=Ng11500;

 always  @(posedge PCLK)
	Ng364<=Ng357;

 always  @(posedge PCLK)
	Ng365<=Ng11501;

 always  @(posedge PCLK)
	Ng366<=Ng365;

 always  @(posedge PCLK)
	Ng367<=Ng11502;

 always  @(posedge PCLK)
	Ng368<=Ng367;

 always  @(posedge PCLK)
	Ng372<=Ng11503;

 always  @(posedge PCLK)
	Ng379<=Ng372;

 always  @(posedge PCLK)
	Ng380<=Ng11504;

 always  @(posedge PCLK)
	Ng381<=Ng380;

 always  @(posedge PCLK)
	Ng382<=Ng11505;

 always  @(posedge PCLK)
	Ng383<=Ng382;

 always  @(posedge PCLK)
	Ng387<=Ng11506;

 always  @(posedge PCLK)
	Ng394<=Ng387;

 always  @(posedge PCLK)
	Ng395<=Ng11507;

 always  @(posedge PCLK)
	Ng396<=Ng395;

 always  @(posedge PCLK)
	Ng397<=Ng11508;

 always  @(posedge PCLK)
	Ng324<=Ng397;

 always  @(posedge PCLK)
	Ng554<=Ng23160;

 always  @(posedge PCLK)
	Ng557<=Ng20556;

 always  @(posedge PCLK)
	Ng510<=Ng20557;

 always  @(posedge PCLK)
	Ng513<=Ng16467;

 always  @(posedge PCLK)
	Ng523<=Ng513;

 always  @(posedge PCLK)
	Ng524<=Ng523;

 always  @(posedge PCLK)
	Ng564<=Ng11512;

 always  @(posedge PCLK)
	Ng569<=Ng564;

 always  @(posedge PCLK)
	Ng570<=Ng11515;

 always  @(posedge PCLK)
	Ng571<=Ng570;

 always  @(posedge PCLK)
	Ng572<=Ng11516;

 always  @(posedge PCLK)
	Ng573<=Ng572;

 always  @(posedge PCLK)
	Ng574<=Ng11517;

 always  @(posedge PCLK)
	Ng565<=Ng574;

 always  @(posedge PCLK)
	Ng566<=Ng11513;

 always  @(posedge PCLK)
	Ng567<=Ng566;

 always  @(posedge PCLK)
	Ng568<=Ng11514;

 always  @(posedge PCLK)
	Ng489<=Ng568;

 always  @(posedge PCLK)
	Ng486<=Ng24292;

 always  @(posedge PCLK)
	Ng487<=Ng24293;

 always  @(posedge PCLK)
	Ng488<=Ng24294;

 always  @(posedge PCLK)
	Ng11512<=Ng25139;

 always  @(posedge PCLK)
	Ng11515<=Ng25131;

 always  @(posedge PCLK)
	Ng11516<=Ng25132;

 always  @(posedge PCLK)
	Ng477<=Ng25136;

 always  @(posedge PCLK)
	Ng478<=Ng25137;

 always  @(posedge PCLK)
	Ng479<=Ng25138;

 always  @(posedge PCLK)
	Ng480<=Ng24289;

 always  @(posedge PCLK)
	Ng484<=Ng24290;

 always  @(posedge PCLK)
	Ng464<=Ng24291;

 always  @(posedge PCLK)
	Ng11517<=Ng25133;

 always  @(posedge PCLK)
	Ng11513<=Ng25134;

 always  @(posedge PCLK)
	Ng11514<=Ng25135;

 always  @(posedge PCLK)
	Ng528<=Ng16468;

 always  @(posedge PCLK)
	Ng535<=Ng528;

 always  @(posedge PCLK)
	Ng542<=Ng535;

 always  @(posedge PCLK)
	Ng543<=Ng19021;

 always  @(posedge PCLK)
	Ng544<=Ng543;

 always  @(posedge PCLK)
	Ng548<=Ng23159;

 always  @(posedge PCLK)
	Ng549<=Ng19022;

 always  @(posedge PCLK)
	Ng8284<=Ng549;

 always  @(posedge PCLK)
	Ng558<=Ng19023;

 always  @(posedge PCLK)
	Ng559<=Ng558;

 always  @(posedge PCLK)
	Ng576<=Ng28219;

 always  @(posedge PCLK)
	Ng577<=Ng28220;

 always  @(posedge PCLK)
	Ng575<=Ng28221;

 always  @(posedge PCLK)
	Ng579<=Ng28222;

 always  @(posedge PCLK)
	Ng580<=Ng28223;

 always  @(posedge PCLK)
	Ng578<=Ng28224;

 always  @(posedge PCLK)
	Ng582<=Ng28225;

 always  @(posedge PCLK)
	Ng583<=Ng28226;

 always  @(posedge PCLK)
	Ng581<=Ng28227;

 always  @(posedge PCLK)
	Ng585<=Ng28228;

 always  @(posedge PCLK)
	Ng586<=Ng28229;

 always  @(posedge PCLK)
	Ng584<=Ng28230;

 always  @(posedge PCLK)
	Ng587<=Ng25985;

 always  @(posedge PCLK)
	Ng590<=Ng25986;

 always  @(posedge PCLK)
	Ng593<=Ng25987;

 always  @(posedge PCLK)
	Ng596<=Ng25988;

 always  @(posedge PCLK)
	Ng599<=Ng25989;

 always  @(posedge PCLK)
	Ng602<=Ng25990;

 always  @(posedge PCLK)
	Ng614<=Ng29135;

 always  @(posedge PCLK)
	Ng617<=Ng29136;

 always  @(posedge PCLK)
	Ng620<=Ng29137;

 always  @(posedge PCLK)
	Ng605<=Ng29132;

 always  @(posedge PCLK)
	Ng608<=Ng29133;

 always  @(posedge PCLK)
	Ng611<=Ng29134;

 always  @(posedge PCLK)
	Ng490<=Ng27194;

 always  @(posedge PCLK)
	Ng493<=Ng27195;

 always  @(posedge PCLK)
	Ng496<=Ng27196;

 always  @(posedge PCLK)
	Ng506<=Ng8284;

 always  @(posedge PCLK)
	Ng507<=Ng24295;

 always  @(posedge PCLK)
	Pg16297<=Ng23154;

 always  @(posedge PCLK)
	Ng525<=Pg16297;

 always  @(posedge PCLK)
	Ng529<=Ng13410;

 always  @(posedge PCLK)
	Ng530<=Ng13411;

 always  @(posedge PCLK)
	Ng531<=Ng13412;

 always  @(posedge PCLK)
	Ng532<=Ng13413;

 always  @(posedge PCLK)
	Ng533<=Ng13414;

 always  @(posedge PCLK)
	Ng534<=Ng13415;

 always  @(posedge PCLK)
	Ng536<=Ng13416;

 always  @(posedge PCLK)
	Ng537<=Ng13417;

 always  @(posedge PCLK)
	Ng538<=Ng25984;

 always  @(posedge PCLK)
	Ng541<=Ng13418;

 always  @(posedge PCLK)
	Ng630<=Ng20558;

 always  @(posedge PCLK)
	Ng659<=Ng21943;

 always  @(posedge PCLK)
	Ng640<=Ng23161;

 always  @(posedge PCLK)
	Ng633<=Ng24296;

 always  @(posedge PCLK)
	Ng653<=Ng25140;

 always  @(posedge PCLK)
	Ng646<=Ng25991;

 always  @(posedge PCLK)
	Ng660<=Ng26691;

 always  @(posedge PCLK)
	Ng672<=Ng27197;

 always  @(posedge PCLK)
	Ng666<=Ng27690;

 always  @(posedge PCLK)
	Ng679<=Ng28231;

 always  @(posedge PCLK)
	Ng686<=Ng28677;

 always  @(posedge PCLK)
	Ng692<=Ng29138;

 always  @(posedge PCLK)
	Ng699<=Ng23162;

 always  @(posedge PCLK)
	Ng700<=Ng23163;

 always  @(posedge PCLK)
	Ng698<=Ng23164;

 always  @(posedge PCLK)
	Ng702<=Ng23165;

 always  @(posedge PCLK)
	Ng703<=Ng23166;

 always  @(posedge PCLK)
	Ng701<=Ng23167;

 always  @(posedge PCLK)
	Ng705<=Ng23168;

 always  @(posedge PCLK)
	Ng706<=Ng23169;

 always  @(posedge PCLK)
	Ng704<=Ng23170;

 always  @(posedge PCLK)
	Ng708<=Ng23171;

 always  @(posedge PCLK)
	Ng709<=Ng23172;

 always  @(posedge PCLK)
	Ng707<=Ng23173;

 always  @(posedge PCLK)
	Ng711<=Ng23174;

 always  @(posedge PCLK)
	Ng712<=Ng23175;

 always  @(posedge PCLK)
	Ng710<=Ng23176;

 always  @(posedge PCLK)
	Ng714<=Ng23177;

 always  @(posedge PCLK)
	Ng715<=Ng23178;

 always  @(posedge PCLK)
	Ng713<=Ng23179;

 always  @(posedge PCLK)
	Ng717<=Ng23180;

 always  @(posedge PCLK)
	Ng718<=Ng23181;

 always  @(posedge PCLK)
	Ng716<=Ng23182;

 always  @(posedge PCLK)
	Ng720<=Ng23183;

 always  @(posedge PCLK)
	Ng721<=Ng23184;

 always  @(posedge PCLK)
	Ng719<=Ng23185;

 always  @(posedge PCLK)
	Ng723<=Ng23186;

 always  @(posedge PCLK)
	Ng724<=Ng23187;

 always  @(posedge PCLK)
	Ng722<=Ng23188;

 always  @(posedge PCLK)
	Ng726<=Ng23189;

 always  @(posedge PCLK)
	Ng727<=Ng23190;

 always  @(posedge PCLK)
	Ng725<=Ng23191;

 always  @(posedge PCLK)
	Ng729<=Ng23192;

 always  @(posedge PCLK)
	Ng730<=Ng23193;

 always  @(posedge PCLK)
	Ng728<=Ng23194;

 always  @(posedge PCLK)
	Ng732<=Ng23195;

 always  @(posedge PCLK)
	Ng733<=Ng23196;

 always  @(posedge PCLK)
	Ng731<=Ng23197;

 always  @(posedge PCLK)
	Ng735<=Ng26692;

 always  @(posedge PCLK)
	Ng736<=Ng26693;

 always  @(posedge PCLK)
	Ng734<=Ng26694;

 always  @(posedge PCLK)
	Ng738<=Ng24297;

 always  @(posedge PCLK)
	Ng739<=Ng24298;

 always  @(posedge PCLK)
	Ng737<=Ng24299;

 always  @(posedge PCLK)
	wire1612<=Ng13457;

 always  @(posedge PCLK)
	wire1594<=wire1612;

 always  @(posedge PCLK)
	Ng853<=wire1594;

 always  @(posedge PCLK)
	Ng818<=Ng24300;

 always  @(posedge PCLK)
	Ng819<=Ng24301;

 always  @(posedge PCLK)
	Ng817<=Ng24302;

 always  @(posedge PCLK)
	Ng821<=Ng24303;

 always  @(posedge PCLK)
	Ng822<=Ng24304;

 always  @(posedge PCLK)
	Ng820<=Ng24305;

 always  @(posedge PCLK)
	Ng830<=Ng24306;

 always  @(posedge PCLK)
	Ng831<=Ng24307;

 always  @(posedge PCLK)
	Ng829<=Ng24308;

 always  @(posedge PCLK)
	Ng833<=Ng24309;

 always  @(posedge PCLK)
	Ng834<=Ng24310;

 always  @(posedge PCLK)
	Ng832<=Ng24311;

 always  @(posedge PCLK)
	Ng836<=Ng24312;

 always  @(posedge PCLK)
	Ng837<=Ng24313;

 always  @(posedge PCLK)
	Ng835<=Ng24314;

 always  @(posedge PCLK)
	Ng839<=Ng24315;

 always  @(posedge PCLK)
	Ng840<=Ng24316;

 always  @(posedge PCLK)
	Ng838<=Ng24317;

 always  @(posedge PCLK)
	Ng842<=Ng24318;

 always  @(posedge PCLK)
	Ng843<=Ng24319;

 always  @(posedge PCLK)
	Ng841<=Ng24320;

 always  @(posedge PCLK)
	Ng845<=Ng24321;

 always  @(posedge PCLK)
	Ng846<=Ng24322;

 always  @(posedge PCLK)
	Ng844<=Ng24323;

 always  @(posedge PCLK)
	Ng848<=Ng24324;

 always  @(posedge PCLK)
	Ng849<=Ng24325;

 always  @(posedge PCLK)
	Ng847<=Ng24326;

 always  @(posedge PCLK)
	Ng851<=Ng24327;

 always  @(posedge PCLK)
	Ng852<=Ng24328;

 always  @(posedge PCLK)
	Ng850<=Ng24329;

 always  @(posedge PCLK)
	Ng857<=Ng26696;

 always  @(posedge PCLK)
	Ng858<=Ng26697;

 always  @(posedge PCLK)
	Ng856<=Ng26698;

 always  @(posedge PCLK)
	Ng860<=Ng26699;

 always  @(posedge PCLK)
	Ng861<=Ng26700;

 always  @(posedge PCLK)
	Ng859<=Ng26701;

 always  @(posedge PCLK)
	Ng863<=Ng26702;

 always  @(posedge PCLK)
	Ng864<=Ng26703;

 always  @(posedge PCLK)
	Ng862<=Ng26704;

 always  @(posedge PCLK)
	Ng866<=Ng26705;

 always  @(posedge PCLK)
	Ng867<=Ng26706;

 always  @(posedge PCLK)
	Ng865<=Ng26707;

 always  @(posedge PCLK)
	Ng873<=Ng30521;

 always  @(posedge PCLK)
	Ng876<=Ng30522;

 always  @(posedge PCLK)
	Ng879<=Ng30523;

 always  @(posedge PCLK)
	Ng918<=Ng30860;

 always  @(posedge PCLK)
	Ng921<=Ng30861;

 always  @(posedge PCLK)
	Ng924<=Ng30862;

 always  @(posedge PCLK)
	Ng882<=Ng30854;

 always  @(posedge PCLK)
	Ng885<=Ng30855;

 always  @(posedge PCLK)
	Ng888<=Ng30856;

 always  @(posedge PCLK)
	Ng927<=Ng30863;

 always  @(posedge PCLK)
	Ng930<=Ng30864;

 always  @(posedge PCLK)
	Ng933<=Ng30865;

 always  @(posedge PCLK)
	Ng891<=Ng30524;

 always  @(posedge PCLK)
	Ng894<=Ng30525;

 always  @(posedge PCLK)
	Ng897<=Ng30526;

 always  @(posedge PCLK)
	Ng936<=Ng30530;

 always  @(posedge PCLK)
	Ng939<=Ng30531;

 always  @(posedge PCLK)
	Ng942<=Ng30532;

 always  @(posedge PCLK)
	Ng900<=Ng30527;

 always  @(posedge PCLK)
	Ng903<=Ng30528;

 always  @(posedge PCLK)
	Ng906<=Ng30529;

 always  @(posedge PCLK)
	Ng945<=Ng30533;

 always  @(posedge PCLK)
	Ng948<=Ng30534;

 always  @(posedge PCLK)
	Ng951<=Ng30535;

 always  @(posedge PCLK)
	Ng909<=Ng30857;

 always  @(posedge PCLK)
	Ng912<=Ng30858;

 always  @(posedge PCLK)
	Ng915<=Ng30859;

 always  @(posedge PCLK)
	Ng954<=Ng30866;

 always  @(posedge PCLK)
	Ng957<=Ng30867;

 always  @(posedge PCLK)
	Ng960<=Ng30868;

 always  @(posedge PCLK)
	Ng780<=Ng25992;

 always  @(posedge PCLK)
	Ng776<=Ng26695;

 always  @(posedge PCLK)
	Ng771<=Ng27198;

 always  @(posedge PCLK)
	Ng767<=Ng27691;

 always  @(posedge PCLK)
	Ng762<=Ng28232;

 always  @(posedge PCLK)
	Ng758<=Ng28678;

 always  @(posedge PCLK)
	Ng753<=Ng29139;

 always  @(posedge PCLK)
	Ng749<=Ng29420;

 always  @(posedge PCLK)
	Ng744<=Ng29634;

 always  @(posedge PCLK)
	Ng740<=Ng29798;

 always  @(posedge PCLK)
	Ng11524<=Ng28233;

 always  @(posedge PCLK)
	Ng11525<=Ng28234;

 always  @(posedge PCLK)
	Ng11526<=Ng28235;

 always  @(posedge PCLK)
	Ng11527<=Ng28236;

 always  @(posedge PCLK)
	Ng11528<=Ng28237;

 always  @(posedge PCLK)
	Ng11529<=Ng28238;

 always  @(posedge PCLK)
	Ng11530<=Ng28239;

 always  @(posedge PCLK)
	Ng11531<=Ng28240;

 always  @(posedge PCLK)
	Ng11532<=Ng28241;

 always  @(posedge PCLK)
	Ng11533<=Ng28242;

 always  @(posedge PCLK)
	Ng11534<=Ng28243;

 always  @(posedge PCLK)
	Ng11535<=Ng28244;

 always  @(posedge PCLK)
	Ng1095<=Ng29421;

 always  @(posedge PCLK)
	Ng1098<=Ng29422;

 always  @(posedge PCLK)
	Ng1101<=Ng29423;

 always  @(posedge PCLK)
	Ng1104<=Ng29638;

 always  @(posedge PCLK)
	Ng1107<=Ng29639;

 always  @(posedge PCLK)
	Ng1110<=Ng29640;

 always  @(posedge PCLK)
	Ng1114<=Ng29424;

 always  @(posedge PCLK)
	Ng1115<=Ng29425;

 always  @(posedge PCLK)
	Ng1113<=Ng29426;

 always  @(posedge PCLK)
	Ng1116<=Ng27692;

 always  @(posedge PCLK)
	Ng1119<=Ng27693;

 always  @(posedge PCLK)
	Ng1122<=Ng27694;

 always  @(posedge PCLK)
	Ng1125<=Ng27695;

 always  @(posedge PCLK)
	Ng1128<=Ng27696;

 always  @(posedge PCLK)
	Ng1131<=Ng27697;

 always  @(posedge PCLK)
	Ng1135<=Ng28679;

 always  @(posedge PCLK)
	Ng1136<=Ng28680;

 always  @(posedge PCLK)
	Ng1134<=Ng28681;

 always  @(posedge PCLK)
	Ng999<=Ng29799;

 always  @(posedge PCLK)
	Ng1000<=Ng29800;

 always  @(posedge PCLK)
	Ng1001<=Ng29801;

 always  @(posedge PCLK)
	Ng1002<=Ng30869;

 always  @(posedge PCLK)
	Ng1003<=Ng30870;

 always  @(posedge PCLK)
	Ng1004<=Ng30871;

 always  @(posedge PCLK)
	Ng1005<=Ng30713;

 always  @(posedge PCLK)
	Ng1006<=Ng30714;

 always  @(posedge PCLK)
	Ng1007<=Ng30715;

 always  @(posedge PCLK)
	Ng1009<=Ng29635;

 always  @(posedge PCLK)
	Ng1010<=Ng29636;

 always  @(posedge PCLK)
	Ng1008<=Ng29637;

 always  @(posedge PCLK)
	Ng1090<=Ng27206;

 always  @(posedge PCLK)
	Ng1091<=Ng27207;

 always  @(posedge PCLK)
	Ng1089<=Ng27208;

 always  @(posedge PCLK)
	Ng1137<=Ng11536;

 always  @(posedge PCLK)
	Ng1138<=Ng1137;

 always  @(posedge PCLK)
	Ng1139<=Ng11537;

 always  @(posedge PCLK)
	Ng1140<=Ng1139;

 always  @(posedge PCLK)
	Ng1141<=Ng11538;

 always  @(posedge PCLK)
	Ng966<=Ng1141;

 always  @(posedge PCLK)
	Ng967<=Ng11518;

 always  @(posedge PCLK)
	Ng968<=Ng967;

 always  @(posedge PCLK)
	Ng969<=Ng11519;

 always  @(posedge PCLK)
	Ng970<=Ng969;

 always  @(posedge PCLK)
	Ng971<=Ng11520;

 always  @(posedge PCLK)
	Ng972<=Ng971;

 always  @(posedge PCLK)
	Ng973<=Ng11521;

 always  @(posedge PCLK)
	Ng974<=Ng973;

 always  @(posedge PCLK)
	Ng975<=Ng11522;

 always  @(posedge PCLK)
	Ng976<=Ng975;

 always  @(posedge PCLK)
	Ng977<=Ng13423;

 always  @(posedge PCLK)
	Ng978<=Ng977;

 always  @(posedge PCLK)
	Ng986<=Ng19024;

 always  @(posedge PCLK)
	Ng992<=Ng27200;

 always  @(posedge PCLK)
	Ng985<=Ng27199;

 always  @(posedge PCLK)
	Ng1029<=Ng11524;

 always  @(posedge PCLK)
	Ng1036<=Ng1029;

 always  @(posedge PCLK)
	Ng1037<=Ng11525;

 always  @(posedge PCLK)
	Ng1038<=Ng1037;

 always  @(posedge PCLK)
	Ng1039<=Ng11526;

 always  @(posedge PCLK)
	Ng1040<=Ng1039;

 always  @(posedge PCLK)
	Ng1044<=Ng11527;

 always  @(posedge PCLK)
	Ng1051<=Ng1044;

 always  @(posedge PCLK)
	Ng1052<=Ng11528;

 always  @(posedge PCLK)
	Ng1053<=Ng1052;

 always  @(posedge PCLK)
	Ng1054<=Ng11529;

 always  @(posedge PCLK)
	Ng1055<=Ng1054;

 always  @(posedge PCLK)
	Ng1059<=Ng11530;

 always  @(posedge PCLK)
	Ng1066<=Ng1059;

 always  @(posedge PCLK)
	Ng1067<=Ng11531;

 always  @(posedge PCLK)
	Ng1068<=Ng1067;

 always  @(posedge PCLK)
	Ng1069<=Ng11532;

 always  @(posedge PCLK)
	Ng1070<=Ng1069;

 always  @(posedge PCLK)
	Ng1074<=Ng11533;

 always  @(posedge PCLK)
	Ng1081<=Ng1074;

 always  @(posedge PCLK)
	Ng1082<=Ng11534;

 always  @(posedge PCLK)
	Ng1083<=Ng1082;

 always  @(posedge PCLK)
	Ng1084<=Ng11535;

 always  @(posedge PCLK)
	Ng1011<=Ng1084;

 always  @(posedge PCLK)
	Ng1240<=Ng23198;

 always  @(posedge PCLK)
	Ng1243<=Ng20560;

 always  @(posedge PCLK)
	Ng1196<=Ng20561;

 always  @(posedge PCLK)
	Ng1199<=Ng16469;

 always  @(posedge PCLK)
	Ng1209<=Ng1199;

 always  @(posedge PCLK)
	Ng1210<=Ng1209;

 always  @(posedge PCLK)
	Ng1250<=Ng11539;

 always  @(posedge PCLK)
	Ng1255<=Ng1250;

 always  @(posedge PCLK)
	Ng1256<=Ng11542;

 always  @(posedge PCLK)
	Ng1257<=Ng1256;

 always  @(posedge PCLK)
	Ng1258<=Ng11543;

 always  @(posedge PCLK)
	Ng1259<=Ng1258;

 always  @(posedge PCLK)
	Ng1260<=Ng11544;

 always  @(posedge PCLK)
	Ng1251<=Ng1260;

 always  @(posedge PCLK)
	Ng1252<=Ng11540;

 always  @(posedge PCLK)
	Ng1253<=Ng1252;

 always  @(posedge PCLK)
	Ng1254<=Ng11541;

 always  @(posedge PCLK)
	Ng1176<=Ng1254;

 always  @(posedge PCLK)
	Ng1173<=Ng24333;

 always  @(posedge PCLK)
	Ng1174<=Ng24334;

 always  @(posedge PCLK)
	Ng1175<=Ng24335;

 always  @(posedge PCLK)
	Ng11539<=Ng25150;

 always  @(posedge PCLK)
	Ng11542<=Ng25142;

 always  @(posedge PCLK)
	Ng11543<=Ng25143;

 always  @(posedge PCLK)
	Ng1164<=Ng25147;

 always  @(posedge PCLK)
	Ng1165<=Ng25148;

 always  @(posedge PCLK)
	Ng1166<=Ng25149;

 always  @(posedge PCLK)
	Ng1167<=Ng24330;

 always  @(posedge PCLK)
	Ng1171<=Ng24331;

 always  @(posedge PCLK)
	Ng1151<=Ng24332;

 always  @(posedge PCLK)
	Ng11544<=Ng25144;

 always  @(posedge PCLK)
	Ng11540<=Ng25145;

 always  @(posedge PCLK)
	Ng11541<=Ng25146;

 always  @(posedge PCLK)
	Ng1214<=Ng16470;

 always  @(posedge PCLK)
	Ng1221<=Ng1214;

 always  @(posedge PCLK)
	Ng1228<=Ng1221;

 always  @(posedge PCLK)
	Ng1229<=Ng19033;

 always  @(posedge PCLK)
	Ng1230<=Ng1229;

 always  @(posedge PCLK)
	Ng1234<=Ng27217;

 always  @(posedge PCLK)
	Ng1235<=Ng19034;

 always  @(posedge PCLK)
	Ng8293<=Ng1235;

 always  @(posedge PCLK)
	Ng1244<=Ng19035;

 always  @(posedge PCLK)
	Ng1245<=Ng1244;

 always  @(posedge PCLK)
	Ng1262<=Ng28245;

 always  @(posedge PCLK)
	Ng1263<=Ng28246;

 always  @(posedge PCLK)
	Ng1261<=Ng28247;

 always  @(posedge PCLK)
	Ng1265<=Ng28248;

 always  @(posedge PCLK)
	Ng1266<=Ng28249;

 always  @(posedge PCLK)
	Ng1264<=Ng28250;

 always  @(posedge PCLK)
	Ng1268<=Ng28251;

 always  @(posedge PCLK)
	Ng1269<=Ng28252;

 always  @(posedge PCLK)
	Ng1267<=Ng28253;

 always  @(posedge PCLK)
	Ng1271<=Ng28254;

 always  @(posedge PCLK)
	Ng1272<=Ng28255;

 always  @(posedge PCLK)
	Ng1270<=Ng28256;

 always  @(posedge PCLK)
	Ng1273<=Ng25994;

 always  @(posedge PCLK)
	Ng1276<=Ng25995;

 always  @(posedge PCLK)
	Ng1279<=Ng25996;

 always  @(posedge PCLK)
	Ng1282<=Ng25997;

 always  @(posedge PCLK)
	Ng1285<=Ng25998;

 always  @(posedge PCLK)
	Ng1288<=Ng25999;

 always  @(posedge PCLK)
	Ng1300<=Ng29143;

 always  @(posedge PCLK)
	Ng1303<=Ng29144;

 always  @(posedge PCLK)
	Ng1306<=Ng29145;

 always  @(posedge PCLK)
	Ng1291<=Ng29140;

 always  @(posedge PCLK)
	Ng1294<=Ng29141;

 always  @(posedge PCLK)
	Ng1297<=Ng29142;

 always  @(posedge PCLK)
	Ng1177<=Ng27209;

 always  @(posedge PCLK)
	Ng1180<=Ng27210;

 always  @(posedge PCLK)
	Ng1183<=Ng27211;

 always  @(posedge PCLK)
	Ng1192<=Ng8293;

 always  @(posedge PCLK)
	Ng1193<=Ng24336;

 always  @(posedge PCLK)
	Pg16355<=Ng27212;

 always  @(posedge PCLK)
	Ng1211<=Pg16355;

 always  @(posedge PCLK)
	Ng1215<=Ng13426;

 always  @(posedge PCLK)
	Ng1216<=Ng13427;

 always  @(posedge PCLK)
	Ng1217<=Ng13428;

 always  @(posedge PCLK)
	Ng1218<=Ng13429;

 always  @(posedge PCLK)
	Ng1219<=Ng13430;

 always  @(posedge PCLK)
	Ng1220<=Ng13431;

 always  @(posedge PCLK)
	Ng1222<=Ng13432;

 always  @(posedge PCLK)
	Ng1223<=Ng13433;

 always  @(posedge PCLK)
	Ng1224<=Ng25993;

 always  @(posedge PCLK)
	Ng1227<=Ng13434;

 always  @(posedge PCLK)
	wire1605<=Ng13475;

 always  @(posedge PCLK)
	wire1603<=wire1605;

 always  @(posedge PCLK)
	Ng1315<=wire1603;

 always  @(posedge PCLK)
	Ng1316<=Ng20562;

 always  @(posedge PCLK)
	Ng1345<=Ng21944;

 always  @(posedge PCLK)
	Ng1326<=Ng23199;

 always  @(posedge PCLK)
	Ng1319<=Ng24337;

 always  @(posedge PCLK)
	Ng1339<=Ng25151;

 always  @(posedge PCLK)
	Ng1332<=Ng26000;

 always  @(posedge PCLK)
	Ng1346<=Ng26708;

 always  @(posedge PCLK)
	Ng1358<=Ng27218;

 always  @(posedge PCLK)
	Ng1352<=Ng27698;

 always  @(posedge PCLK)
	Ng1365<=Ng28257;

 always  @(posedge PCLK)
	Ng1372<=Ng28682;

 always  @(posedge PCLK)
	Ng1378<=Ng29146;

 always  @(posedge PCLK)
	Ng1385<=Ng23200;

 always  @(posedge PCLK)
	Ng1386<=Ng23201;

 always  @(posedge PCLK)
	Ng1384<=Ng23202;

 always  @(posedge PCLK)
	Ng1388<=Ng23203;

 always  @(posedge PCLK)
	Ng1389<=Ng23204;

 always  @(posedge PCLK)
	Ng1387<=Ng23205;

 always  @(posedge PCLK)
	Ng1391<=Ng23206;

 always  @(posedge PCLK)
	Ng1392<=Ng23207;

 always  @(posedge PCLK)
	Ng1390<=Ng23208;

 always  @(posedge PCLK)
	Ng1394<=Ng23209;

 always  @(posedge PCLK)
	Ng1395<=Ng23210;

 always  @(posedge PCLK)
	Ng1393<=Ng23211;

 always  @(posedge PCLK)
	Ng1397<=Ng23212;

 always  @(posedge PCLK)
	Ng1398<=Ng23213;

 always  @(posedge PCLK)
	Ng1396<=Ng23214;

 always  @(posedge PCLK)
	Ng1400<=Ng23215;

 always  @(posedge PCLK)
	Ng1401<=Ng23216;

 always  @(posedge PCLK)
	Ng1399<=Ng23217;

 always  @(posedge PCLK)
	Ng1403<=Ng23218;

 always  @(posedge PCLK)
	Ng1404<=Ng23219;

 always  @(posedge PCLK)
	Ng1402<=Ng23220;

 always  @(posedge PCLK)
	Ng1406<=Ng23221;

 always  @(posedge PCLK)
	Ng1407<=Ng23222;

 always  @(posedge PCLK)
	Ng1405<=Ng23223;

 always  @(posedge PCLK)
	Ng1409<=Ng23224;

 always  @(posedge PCLK)
	Ng1410<=Ng23225;

 always  @(posedge PCLK)
	Ng1408<=Ng23226;

 always  @(posedge PCLK)
	Ng1412<=Ng23227;

 always  @(posedge PCLK)
	Ng1413<=Ng23228;

 always  @(posedge PCLK)
	Ng1411<=Ng23229;

 always  @(posedge PCLK)
	Ng1415<=Ng23230;

 always  @(posedge PCLK)
	Ng1416<=Ng23231;

 always  @(posedge PCLK)
	Ng1414<=Ng23232;

 always  @(posedge PCLK)
	Ng1418<=Ng23233;

 always  @(posedge PCLK)
	Ng1419<=Ng23234;

 always  @(posedge PCLK)
	Ng1417<=Ng23235;

 always  @(posedge PCLK)
	Ng1421<=Ng26709;

 always  @(posedge PCLK)
	Ng1422<=Ng26710;

 always  @(posedge PCLK)
	Ng1420<=Ng26711;

 always  @(posedge PCLK)
	Ng1424<=Ng24338;

 always  @(posedge PCLK)
	Ng1425<=Ng24339;

 always  @(posedge PCLK)
	Ng1423<=Ng24340;

 always  @(posedge PCLK)
	Ng1512<=Ng24341;

 always  @(posedge PCLK)
	Ng1513<=Ng24342;

 always  @(posedge PCLK)
	Ng1511<=Ng24343;

 always  @(posedge PCLK)
	Ng1515<=Ng24344;

 always  @(posedge PCLK)
	Ng1516<=Ng24345;

 always  @(posedge PCLK)
	Ng1514<=Ng24346;

 always  @(posedge PCLK)
	Ng1524<=Ng24347;

 always  @(posedge PCLK)
	Ng1525<=Ng24348;

 always  @(posedge PCLK)
	Ng1523<=Ng24349;

 always  @(posedge PCLK)
	Ng1527<=Ng24350;

 always  @(posedge PCLK)
	Ng1528<=Ng24351;

 always  @(posedge PCLK)
	Ng1526<=Ng24352;

 always  @(posedge PCLK)
	Ng1530<=Ng24353;

 always  @(posedge PCLK)
	Ng1531<=Ng24354;

 always  @(posedge PCLK)
	Ng1529<=Ng24355;

 always  @(posedge PCLK)
	Ng1533<=Ng24356;

 always  @(posedge PCLK)
	Ng1534<=Ng24357;

 always  @(posedge PCLK)
	Ng1532<=Ng24358;

 always  @(posedge PCLK)
	Ng1536<=Ng24359;

 always  @(posedge PCLK)
	Ng1537<=Ng24360;

 always  @(posedge PCLK)
	Ng1535<=Ng24361;

 always  @(posedge PCLK)
	Ng1539<=Ng24362;

 always  @(posedge PCLK)
	Ng1540<=Ng24363;

 always  @(posedge PCLK)
	Ng1538<=Ng24364;

 always  @(posedge PCLK)
	Ng1542<=Ng24365;

 always  @(posedge PCLK)
	Ng1543<=Ng24366;

 always  @(posedge PCLK)
	Ng1541<=Ng24367;

 always  @(posedge PCLK)
	Ng1545<=Ng24368;

 always  @(posedge PCLK)
	Ng1546<=Ng24369;

 always  @(posedge PCLK)
	Ng1544<=Ng24370;

 always  @(posedge PCLK)
	Ng1551<=Ng26713;

 always  @(posedge PCLK)
	Ng1552<=Ng26714;

 always  @(posedge PCLK)
	Ng1550<=Ng26715;

 always  @(posedge PCLK)
	Ng1554<=Ng26716;

 always  @(posedge PCLK)
	Ng1555<=Ng26717;

 always  @(posedge PCLK)
	Ng1553<=Ng26718;

 always  @(posedge PCLK)
	Ng1557<=Ng26719;

 always  @(posedge PCLK)
	Ng1558<=Ng26720;

 always  @(posedge PCLK)
	Ng1556<=Ng26721;

 always  @(posedge PCLK)
	Ng1560<=Ng26722;

 always  @(posedge PCLK)
	Ng1561<=Ng26723;

 always  @(posedge PCLK)
	Ng1559<=Ng26724;

 always  @(posedge PCLK)
	Ng1567<=Ng30536;

 always  @(posedge PCLK)
	Ng1570<=Ng30537;

 always  @(posedge PCLK)
	Ng1573<=Ng30538;

 always  @(posedge PCLK)
	Ng1612<=Ng30878;

 always  @(posedge PCLK)
	Ng1615<=Ng30879;

 always  @(posedge PCLK)
	Ng1618<=Ng30880;

 always  @(posedge PCLK)
	Ng1576<=Ng30872;

 always  @(posedge PCLK)
	Ng1579<=Ng30873;

 always  @(posedge PCLK)
	Ng1582<=Ng30874;

 always  @(posedge PCLK)
	Ng1621<=Ng30881;

 always  @(posedge PCLK)
	Ng1624<=Ng30882;

 always  @(posedge PCLK)
	Ng1627<=Ng30883;

 always  @(posedge PCLK)
	Ng1585<=Ng30539;

 always  @(posedge PCLK)
	Ng1588<=Ng30540;

 always  @(posedge PCLK)
	Ng1591<=Ng30541;

 always  @(posedge PCLK)
	Ng1630<=Ng30545;

 always  @(posedge PCLK)
	Ng1633<=Ng30546;

 always  @(posedge PCLK)
	Ng1636<=Ng30547;

 always  @(posedge PCLK)
	Ng1594<=Ng30542;

 always  @(posedge PCLK)
	Ng1597<=Ng30543;

 always  @(posedge PCLK)
	Ng1600<=Ng30544;

 always  @(posedge PCLK)
	Ng1639<=Ng30548;

 always  @(posedge PCLK)
	Ng1642<=Ng30549;

 always  @(posedge PCLK)
	Ng1645<=Ng30550;

 always  @(posedge PCLK)
	Ng1603<=Ng30875;

 always  @(posedge PCLK)
	Ng1606<=Ng30876;

 always  @(posedge PCLK)
	Ng1609<=Ng30877;

 always  @(posedge PCLK)
	Ng1648<=Ng30884;

 always  @(posedge PCLK)
	Ng1651<=Ng30885;

 always  @(posedge PCLK)
	Ng1654<=Ng30886;

 always  @(posedge PCLK)
	Ng1466<=Ng26001;

 always  @(posedge PCLK)
	Ng1462<=Ng26712;

 always  @(posedge PCLK)
	Ng1457<=Ng27219;

 always  @(posedge PCLK)
	Ng1453<=Ng27699;

 always  @(posedge PCLK)
	Ng1448<=Ng28258;

 always  @(posedge PCLK)
	Ng1444<=Ng28683;

 always  @(posedge PCLK)
	Ng1439<=Ng29147;

 always  @(posedge PCLK)
	Ng1435<=Ng29427;

 always  @(posedge PCLK)
	Ng1430<=Ng29641;

 always  @(posedge PCLK)
	Ng1426<=Ng29802;

 always  @(posedge PCLK)
	Ng11551<=Ng28259;

 always  @(posedge PCLK)
	Ng11552<=Ng28260;

 always  @(posedge PCLK)
	Ng11553<=Ng28261;

 always  @(posedge PCLK)
	Ng11554<=Ng28262;

 always  @(posedge PCLK)
	Ng11555<=Ng28263;

 always  @(posedge PCLK)
	Ng11556<=Ng28264;

 always  @(posedge PCLK)
	Ng11557<=Ng28265;

 always  @(posedge PCLK)
	Ng11558<=Ng28266;

 always  @(posedge PCLK)
	Ng11559<=Ng28267;

 always  @(posedge PCLK)
	Ng11560<=Ng28268;

 always  @(posedge PCLK)
	Ng11561<=Ng28269;

 always  @(posedge PCLK)
	Ng11562<=Ng28270;

 always  @(posedge PCLK)
	Ng1789<=Ng29434;

 always  @(posedge PCLK)
	Ng1792<=Ng29435;

 always  @(posedge PCLK)
	Ng1795<=Ng29436;

 always  @(posedge PCLK)
	Ng1798<=Ng29645;

 always  @(posedge PCLK)
	Ng1801<=Ng29646;

 always  @(posedge PCLK)
	Ng1804<=Ng29647;

 always  @(posedge PCLK)
	Ng1808<=Ng29437;

 always  @(posedge PCLK)
	Ng1809<=Ng29438;

 always  @(posedge PCLK)
	Ng1807<=Ng29439;

 always  @(posedge PCLK)
	Ng1810<=Ng27700;

 always  @(posedge PCLK)
	Ng1813<=Ng27701;

 always  @(posedge PCLK)
	Ng1816<=Ng27702;

 always  @(posedge PCLK)
	Ng1819<=Ng27703;

 always  @(posedge PCLK)
	Ng1822<=Ng27704;

 always  @(posedge PCLK)
	Ng1825<=Ng27705;

 always  @(posedge PCLK)
	Ng1829<=Ng28684;

 always  @(posedge PCLK)
	Ng1830<=Ng28685;

 always  @(posedge PCLK)
	Ng1828<=Ng28686;

 always  @(posedge PCLK)
	Ng1693<=Ng29803;

 always  @(posedge PCLK)
	Ng1694<=Ng29804;

 always  @(posedge PCLK)
	Ng1695<=Ng29805;

 always  @(posedge PCLK)
	Ng1696<=Ng30887;

 always  @(posedge PCLK)
	Ng1697<=Ng30888;

 always  @(posedge PCLK)
	Ng1698<=Ng30889;

 always  @(posedge PCLK)
	Ng1699<=Ng30716;

 always  @(posedge PCLK)
	Ng1700<=Ng30717;

 always  @(posedge PCLK)
	Ng1701<=Ng30718;

 always  @(posedge PCLK)
	Ng1703<=Ng29642;

 always  @(posedge PCLK)
	Ng1704<=Ng29643;

 always  @(posedge PCLK)
	Ng1702<=Ng29644;

 always  @(posedge PCLK)
	Ng1784<=Ng27221;

 always  @(posedge PCLK)
	Ng1785<=Ng27222;

 always  @(posedge PCLK)
	Ng1783<=Ng27223;

 always  @(posedge PCLK)
	Ng1831<=Ng11563;

 always  @(posedge PCLK)
	Ng1832<=Ng1831;

 always  @(posedge PCLK)
	Ng1833<=Ng11564;

 always  @(posedge PCLK)
	Ng1834<=Ng1833;

 always  @(posedge PCLK)
	Ng1835<=Ng11565;

 always  @(posedge PCLK)
	Ng1660<=Ng1835;

 always  @(posedge PCLK)
	Ng1661<=Ng11545;

 always  @(posedge PCLK)
	Ng1662<=Ng1661;

 always  @(posedge PCLK)
	Ng1663<=Ng11546;

 always  @(posedge PCLK)
	Ng1664<=Ng1663;

 always  @(posedge PCLK)
	Ng1665<=Ng11547;

 always  @(posedge PCLK)
	Ng1666<=Ng1665;

 always  @(posedge PCLK)
	Ng1667<=Ng11548;

 always  @(posedge PCLK)
	Ng1668<=Ng1667;

 always  @(posedge PCLK)
	Ng1669<=Ng11549;

 always  @(posedge PCLK)
	Ng1670<=Ng1669;

 always  @(posedge PCLK)
	Ng1671<=Ng13439;

 always  @(posedge PCLK)
	Ng1672<=Ng1671;

 always  @(posedge PCLK)
	Ng1680<=Ng19036;

 always  @(posedge PCLK)
	Ng1686<=Ng29428;

 always  @(posedge PCLK)
	Ng1679<=Ng27220;

 always  @(posedge PCLK)
	Ng1723<=Ng11551;

 always  @(posedge PCLK)
	Ng1730<=Ng1723;

 always  @(posedge PCLK)
	Ng1731<=Ng11552;

 always  @(posedge PCLK)
	Ng1732<=Ng1731;

 always  @(posedge PCLK)
	Ng1733<=Ng11553;

 always  @(posedge PCLK)
	Ng1734<=Ng1733;

 always  @(posedge PCLK)
	Ng1738<=Ng11554;

 always  @(posedge PCLK)
	Ng1745<=Ng1738;

 always  @(posedge PCLK)
	Ng1746<=Ng11555;

 always  @(posedge PCLK)
	Ng1747<=Ng1746;

 always  @(posedge PCLK)
	Ng1748<=Ng11556;

 always  @(posedge PCLK)
	Ng1749<=Ng1748;

 always  @(posedge PCLK)
	Ng1753<=Ng11557;

 always  @(posedge PCLK)
	Ng1760<=Ng1753;

 always  @(posedge PCLK)
	Ng1761<=Ng11558;

 always  @(posedge PCLK)
	Ng1762<=Ng1761;

 always  @(posedge PCLK)
	Ng1763<=Ng11559;

 always  @(posedge PCLK)
	Ng1764<=Ng1763;

 always  @(posedge PCLK)
	Ng1768<=Ng11560;

 always  @(posedge PCLK)
	Ng1775<=Ng1768;

 always  @(posedge PCLK)
	Ng1776<=Ng11561;

 always  @(posedge PCLK)
	Ng1777<=Ng1776;

 always  @(posedge PCLK)
	Ng1778<=Ng11562;

 always  @(posedge PCLK)
	Ng1705<=Ng1778;

 always  @(posedge PCLK)
	Ng1934<=Ng23236;

 always  @(posedge PCLK)
	Ng1937<=Ng20564;

 always  @(posedge PCLK)
	Ng1890<=Ng20565;

 always  @(posedge PCLK)
	Ng1893<=Ng16471;

 always  @(posedge PCLK)
	Ng1903<=Ng1893;

 always  @(posedge PCLK)
	Ng1904<=Ng1903;

 always  @(posedge PCLK)
	Ng1944<=Ng11566;

 always  @(posedge PCLK)
	Ng1949<=Ng1944;

 always  @(posedge PCLK)
	Ng1950<=Ng11569;

 always  @(posedge PCLK)
	Ng1951<=Ng1950;

 always  @(posedge PCLK)
	Ng1952<=Ng11570;

 always  @(posedge PCLK)
	Ng1953<=Ng1952;

 always  @(posedge PCLK)
	Ng1954<=Ng11571;

 always  @(posedge PCLK)
	Ng1945<=Ng1954;

 always  @(posedge PCLK)
	Ng1946<=Ng11567;

 always  @(posedge PCLK)
	Ng1947<=Ng1946;

 always  @(posedge PCLK)
	Ng1948<=Ng11568;

 always  @(posedge PCLK)
	Ng1870<=Ng1948;

 always  @(posedge PCLK)
	Ng1867<=Ng24374;

 always  @(posedge PCLK)
	Ng1868<=Ng24375;

 always  @(posedge PCLK)
	Ng1869<=Ng24376;

 always  @(posedge PCLK)
	Ng11566<=Ng25161;

 always  @(posedge PCLK)
	Ng11569<=Ng25153;

 always  @(posedge PCLK)
	Ng11570<=Ng25154;

 always  @(posedge PCLK)
	Ng1858<=Ng25158;

 always  @(posedge PCLK)
	Ng1859<=Ng25159;

 always  @(posedge PCLK)
	Ng1860<=Ng25160;

 always  @(posedge PCLK)
	Ng1861<=Ng24371;

 always  @(posedge PCLK)
	Ng1865<=Ng24372;

 always  @(posedge PCLK)
	Ng1845<=Ng24373;

 always  @(posedge PCLK)
	Ng11571<=Ng25155;

 always  @(posedge PCLK)
	Ng11567<=Ng25156;

 always  @(posedge PCLK)
	Ng11568<=Ng25157;

 always  @(posedge PCLK)
	Ng1908<=Ng16472;

 always  @(posedge PCLK)
	Ng1915<=Ng1908;

 always  @(posedge PCLK)
	Ng1922<=Ng1915;

 always  @(posedge PCLK)
	Ng1923<=Ng19045;

 always  @(posedge PCLK)
	Ng1924<=Ng1923;

 always  @(posedge PCLK)
	Ng1928<=Ng29445;

 always  @(posedge PCLK)
	Ng1929<=Ng19046;

 always  @(posedge PCLK)
	Ng8302<=Ng1929;

 always  @(posedge PCLK)
	Ng1938<=Ng19047;

 always  @(posedge PCLK)
	Ng1939<=Ng1938;

 always  @(posedge PCLK)
	Ng1956<=Ng28271;

 always  @(posedge PCLK)
	Ng1957<=Ng28272;

 always  @(posedge PCLK)
	Ng1955<=Ng28273;

 always  @(posedge PCLK)
	Ng1959<=Ng28274;

 always  @(posedge PCLK)
	Ng1960<=Ng28275;

 always  @(posedge PCLK)
	Ng1958<=Ng28276;

 always  @(posedge PCLK)
	Ng1962<=Ng28277;

 always  @(posedge PCLK)
	Ng1963<=Ng28278;

 always  @(posedge PCLK)
	Ng1961<=Ng28279;

 always  @(posedge PCLK)
	Ng1965<=Ng28280;

 always  @(posedge PCLK)
	Ng1966<=Ng28281;

 always  @(posedge PCLK)
	Ng1964<=Ng28282;

 always  @(posedge PCLK)
	Ng1967<=Ng26003;

 always  @(posedge PCLK)
	Ng1970<=Ng26004;

 always  @(posedge PCLK)
	Ng1973<=Ng26005;

 always  @(posedge PCLK)
	Ng1976<=Ng26006;

 always  @(posedge PCLK)
	Ng1979<=Ng26007;

 always  @(posedge PCLK)
	Ng1982<=Ng26008;

 always  @(posedge PCLK)
	Ng1994<=Ng29151;

 always  @(posedge PCLK)
	Ng1997<=Ng29152;

 always  @(posedge PCLK)
	Ng2000<=Ng29153;

 always  @(posedge PCLK)
	Ng1985<=Ng29148;

 always  @(posedge PCLK)
	Ng1988<=Ng29149;

 always  @(posedge PCLK)
	Ng1991<=Ng29150;

 always  @(posedge PCLK)
	Ng1871<=Ng27224;

 always  @(posedge PCLK)
	Ng1874<=Ng27225;

 always  @(posedge PCLK)
	Ng1877<=Ng27226;

 always  @(posedge PCLK)
	Ng1886<=Ng8302;

 always  @(posedge PCLK)
	Ng1887<=Ng24377;

 always  @(posedge PCLK)
	Pg16399<=Ng29440;

 always  @(posedge PCLK)
	Ng1905<=Pg16399;

 always  @(posedge PCLK)
	Ng1909<=Ng13442;

 always  @(posedge PCLK)
	Ng1910<=Ng13443;

 always  @(posedge PCLK)
	Ng1911<=Ng13444;

 always  @(posedge PCLK)
	Ng1912<=Ng13445;

 always  @(posedge PCLK)
	Ng1913<=Ng13446;

 always  @(posedge PCLK)
	Ng1914<=Ng13447;

 always  @(posedge PCLK)
	Ng1916<=Ng13448;

 always  @(posedge PCLK)
	Ng1917<=Ng13449;

 always  @(posedge PCLK)
	Ng1918<=Ng26002;

 always  @(posedge PCLK)
	Ng1921<=Ng13450;

 always  @(posedge PCLK)
	Ng2010<=Ng20566;

 always  @(posedge PCLK)
	Ng2039<=Ng21945;

 always  @(posedge PCLK)
	Ng2020<=Ng23237;

 always  @(posedge PCLK)
	Ng2013<=Ng24378;

 always  @(posedge PCLK)
	Ng2033<=Ng25162;

 always  @(posedge PCLK)
	Ng2026<=Ng26009;

 always  @(posedge PCLK)
	Ng2040<=Ng26725;

 always  @(posedge PCLK)
	Ng2052<=Ng27227;

 always  @(posedge PCLK)
	Ng2046<=Ng27706;

 always  @(posedge PCLK)
	Ng2059<=Ng28283;

 always  @(posedge PCLK)
	Ng2066<=Ng28687;

 always  @(posedge PCLK)
	Ng2072<=Ng29154;

 always  @(posedge PCLK)
	Ng2079<=Ng23238;

 always  @(posedge PCLK)
	Ng2080<=Ng23239;

 always  @(posedge PCLK)
	Ng2078<=Ng23240;

 always  @(posedge PCLK)
	Ng2082<=Ng23241;

 always  @(posedge PCLK)
	Ng2083<=Ng23242;

 always  @(posedge PCLK)
	Ng2081<=Ng23243;

 always  @(posedge PCLK)
	Ng2085<=Ng23244;

 always  @(posedge PCLK)
	Ng2086<=Ng23245;

 always  @(posedge PCLK)
	Ng2084<=Ng23246;

 always  @(posedge PCLK)
	Ng2088<=Ng23247;

 always  @(posedge PCLK)
	Ng2089<=Ng23248;

 always  @(posedge PCLK)
	Ng2087<=Ng23249;

 always  @(posedge PCLK)
	Ng2091<=Ng23250;

 always  @(posedge PCLK)
	Ng2092<=Ng23251;

 always  @(posedge PCLK)
	Ng2090<=Ng23252;

 always  @(posedge PCLK)
	Ng2094<=Ng23253;

 always  @(posedge PCLK)
	Ng2095<=Ng23254;

 always  @(posedge PCLK)
	Ng2093<=Ng23255;

 always  @(posedge PCLK)
	Ng2097<=Ng23256;

 always  @(posedge PCLK)
	Ng2098<=Ng23257;

 always  @(posedge PCLK)
	Ng2096<=Ng23258;

 always  @(posedge PCLK)
	Ng2100<=Ng23259;

 always  @(posedge PCLK)
	Ng2101<=Ng23260;

 always  @(posedge PCLK)
	Ng2099<=Ng23261;

 always  @(posedge PCLK)
	Ng2103<=Ng23262;

 always  @(posedge PCLK)
	Ng2104<=Ng23263;

 always  @(posedge PCLK)
	Ng2102<=Ng23264;

 always  @(posedge PCLK)
	Ng2106<=Ng23265;

 always  @(posedge PCLK)
	Ng2107<=Ng23266;

 always  @(posedge PCLK)
	Ng2105<=Ng23267;

 always  @(posedge PCLK)
	Ng2109<=Ng23268;

 always  @(posedge PCLK)
	Ng2110<=Ng23269;

 always  @(posedge PCLK)
	Ng2108<=Ng23270;

 always  @(posedge PCLK)
	Ng2112<=Ng23271;

 always  @(posedge PCLK)
	Ng2113<=Ng23272;

 always  @(posedge PCLK)
	Ng2111<=Ng23273;

 always  @(posedge PCLK)
	Ng2115<=Ng26726;

 always  @(posedge PCLK)
	Ng2116<=Ng26727;

 always  @(posedge PCLK)
	Ng2114<=Ng26728;

 always  @(posedge PCLK)
	Ng2118<=Ng24379;

 always  @(posedge PCLK)
	Ng2119<=Ng24380;

 always  @(posedge PCLK)
	Ng2117<=Ng24381;

 always  @(posedge PCLK)
	Ng2206<=Ng24382;

 always  @(posedge PCLK)
	Ng2207<=Ng24383;

 always  @(posedge PCLK)
	Ng2205<=Ng24384;

 always  @(posedge PCLK)
	Ng2209<=Ng24385;

 always  @(posedge PCLK)
	Ng2210<=Ng24386;

 always  @(posedge PCLK)
	Ng2208<=Ng24387;

 always  @(posedge PCLK)
	Ng2218<=Ng24388;

 always  @(posedge PCLK)
	Ng2219<=Ng24389;

 always  @(posedge PCLK)
	Ng2217<=Ng24390;

 always  @(posedge PCLK)
	Ng2221<=Ng24391;

 always  @(posedge PCLK)
	Ng2222<=Ng24392;

 always  @(posedge PCLK)
	Ng2220<=Ng24393;

 always  @(posedge PCLK)
	Ng2224<=Ng24394;

 always  @(posedge PCLK)
	Ng2225<=Ng24395;

 always  @(posedge PCLK)
	Ng2223<=Ng24396;

 always  @(posedge PCLK)
	Ng2227<=Ng24397;

 always  @(posedge PCLK)
	Ng2228<=Ng24398;

 always  @(posedge PCLK)
	Ng2226<=Ng24399;

 always  @(posedge PCLK)
	Ng2230<=Ng24400;

 always  @(posedge PCLK)
	Ng2231<=Ng24401;

 always  @(posedge PCLK)
	Ng2229<=Ng24402;

 always  @(posedge PCLK)
	Ng2233<=Ng24403;

 always  @(posedge PCLK)
	Ng2234<=Ng24404;

 always  @(posedge PCLK)
	Ng2232<=Ng24405;

 always  @(posedge PCLK)
	Ng2236<=Ng24406;

 always  @(posedge PCLK)
	Ng2237<=Ng24407;

 always  @(posedge PCLK)
	Ng2235<=Ng24408;

 always  @(posedge PCLK)
	Ng2239<=Ng24409;

 always  @(posedge PCLK)
	Ng2240<=Ng24410;

 always  @(posedge PCLK)
	Ng2238<=Ng24411;

 always  @(posedge PCLK)
	Ng2245<=Ng26730;

 always  @(posedge PCLK)
	Ng2246<=Ng26731;

 always  @(posedge PCLK)
	Ng2244<=Ng26732;

 always  @(posedge PCLK)
	Ng2248<=Ng26733;

 always  @(posedge PCLK)
	Ng2249<=Ng26734;

 always  @(posedge PCLK)
	Ng2247<=Ng26735;

 always  @(posedge PCLK)
	Ng2251<=Ng26736;

 always  @(posedge PCLK)
	Ng2252<=Ng26737;

 always  @(posedge PCLK)
	Ng2250<=Ng26738;

 always  @(posedge PCLK)
	Ng2254<=Ng26739;

 always  @(posedge PCLK)
	Ng2255<=Ng26740;

 always  @(posedge PCLK)
	Ng2253<=Ng26741;

 always  @(posedge PCLK)
	Ng2261<=Ng30551;

 always  @(posedge PCLK)
	Ng2264<=Ng30552;

 always  @(posedge PCLK)
	Ng2267<=Ng30553;

 always  @(posedge PCLK)
	Ng2306<=Ng30896;

 always  @(posedge PCLK)
	Ng2309<=Ng30897;

 always  @(posedge PCLK)
	Ng2312<=Ng30898;

 always  @(posedge PCLK)
	Ng2270<=Ng30890;

 always  @(posedge PCLK)
	Ng2273<=Ng30891;

 always  @(posedge PCLK)
	Ng2276<=Ng30892;

 always  @(posedge PCLK)
	Ng2315<=Ng30899;

 always  @(posedge PCLK)
	Ng2318<=Ng30900;

 always  @(posedge PCLK)
	Ng2321<=Ng30901;

 always  @(posedge PCLK)
	Ng2279<=Ng30554;

 always  @(posedge PCLK)
	Ng2282<=Ng30555;

 always  @(posedge PCLK)
	Ng2285<=Ng30556;

 always  @(posedge PCLK)
	Ng2324<=Ng30560;

 always  @(posedge PCLK)
	Ng2327<=Ng30561;

 always  @(posedge PCLK)
	Ng2330<=Ng30562;

 always  @(posedge PCLK)
	Ng2288<=Ng30557;

 always  @(posedge PCLK)
	Ng2291<=Ng30558;

 always  @(posedge PCLK)
	Ng2294<=Ng30559;

 always  @(posedge PCLK)
	Ng2333<=Ng30563;

 always  @(posedge PCLK)
	Ng2336<=Ng30564;

 always  @(posedge PCLK)
	Ng2339<=Ng30565;

 always  @(posedge PCLK)
	Ng2297<=Ng30893;

 always  @(posedge PCLK)
	Ng2300<=Ng30894;

 always  @(posedge PCLK)
	Ng2303<=Ng30895;

 always  @(posedge PCLK)
	Ng2342<=Ng30902;

 always  @(posedge PCLK)
	Ng2345<=Ng30903;

 always  @(posedge PCLK)
	Ng2348<=Ng30904;

 always  @(posedge PCLK)
	Ng2160<=Ng26010;

 always  @(posedge PCLK)
	Ng2156<=Ng26729;

 always  @(posedge PCLK)
	Ng2151<=Ng27228;

 always  @(posedge PCLK)
	Ng2147<=Ng27707;

 always  @(posedge PCLK)
	Ng2142<=Ng28284;

 always  @(posedge PCLK)
	Ng2138<=Ng28688;

 always  @(posedge PCLK)
	Ng2133<=Ng29155;

 always  @(posedge PCLK)
	Ng2129<=Ng29446;

 always  @(posedge PCLK)
	Ng2124<=Ng29648;

 always  @(posedge PCLK)
	Ng2120<=Ng29806;

 always  @(posedge PCLK)
	Ng2256<=Ng20567;

 always  @(posedge PCLK)
	wire1609<=Ng2256;

 always  @(posedge PCLK)
	Ng2257<=wire1609;

 always  @(posedge PCLK)
	Ng11578<=Ng28285;

 always  @(posedge PCLK)
	Ng11579<=Ng28286;

 always  @(posedge PCLK)
	Ng11580<=Ng28287;

 always  @(posedge PCLK)
	Ng11581<=Ng28288;

 always  @(posedge PCLK)
	Ng11582<=Ng28289;

 always  @(posedge PCLK)
	Ng11583<=Ng28290;

 always  @(posedge PCLK)
	Ng11584<=Ng28291;

 always  @(posedge PCLK)
	Ng11585<=Ng28292;

 always  @(posedge PCLK)
	Ng11586<=Ng28293;

 always  @(posedge PCLK)
	Ng11587<=Ng28294;

 always  @(posedge PCLK)
	Ng11588<=Ng28295;

 always  @(posedge PCLK)
	Ng11589<=Ng28296;

 always  @(posedge PCLK)
	Ng2483<=Ng29447;

 always  @(posedge PCLK)
	Ng2486<=Ng29448;

 always  @(posedge PCLK)
	Ng2489<=Ng29449;

 always  @(posedge PCLK)
	Ng2492<=Ng29652;

 always  @(posedge PCLK)
	Ng2495<=Ng29653;

 always  @(posedge PCLK)
	Ng2498<=Ng29654;

 always  @(posedge PCLK)
	Ng2502<=Ng29450;

 always  @(posedge PCLK)
	Ng2503<=Ng29451;

 always  @(posedge PCLK)
	Ng2501<=Ng29452;

 always  @(posedge PCLK)
	Ng2504<=Ng27708;

 always  @(posedge PCLK)
	Ng2507<=Ng27709;

 always  @(posedge PCLK)
	Ng2510<=Ng27710;

 always  @(posedge PCLK)
	Ng2513<=Ng27711;

 always  @(posedge PCLK)
	Ng2516<=Ng27712;

 always  @(posedge PCLK)
	Ng2519<=Ng27713;

 always  @(posedge PCLK)
	Ng2523<=Ng28689;

 always  @(posedge PCLK)
	Ng2524<=Ng28690;

 always  @(posedge PCLK)
	Ng2522<=Ng28691;

 always  @(posedge PCLK)
	Ng2387<=Ng29807;

 always  @(posedge PCLK)
	Ng2388<=Ng29808;

 always  @(posedge PCLK)
	Ng2389<=Ng29809;

 always  @(posedge PCLK)
	Ng2390<=Ng30905;

 always  @(posedge PCLK)
	Ng2391<=Ng30906;

 always  @(posedge PCLK)
	Ng2392<=Ng30907;

 always  @(posedge PCLK)
	Ng2393<=Ng30719;

 always  @(posedge PCLK)
	Ng2394<=Ng30720;

 always  @(posedge PCLK)
	Ng2395<=Ng30721;

 always  @(posedge PCLK)
	Ng2397<=Ng29649;

 always  @(posedge PCLK)
	Ng2398<=Ng29650;

 always  @(posedge PCLK)
	Ng2396<=Ng29651;

 always  @(posedge PCLK)
	Ng2478<=Ng27230;

 always  @(posedge PCLK)
	Ng2479<=Ng27231;

 always  @(posedge PCLK)
	Ng2477<=Ng27232;

 always  @(posedge PCLK)
	Ng2525<=Ng11590;

 always  @(posedge PCLK)
	Ng2526<=Ng2525;

 always  @(posedge PCLK)
	Ng2527<=Ng11591;

 always  @(posedge PCLK)
	Ng2528<=Ng2527;

 always  @(posedge PCLK)
	Ng2529<=Ng11592;

 always  @(posedge PCLK)
	Ng2354<=Ng2529;

 always  @(posedge PCLK)
	Ng2355<=Ng11572;

 always  @(posedge PCLK)
	Ng2356<=Ng2355;

 always  @(posedge PCLK)
	Ng2357<=Ng11573;

 always  @(posedge PCLK)
	Ng2358<=Ng2357;

 always  @(posedge PCLK)
	Ng2359<=Ng11574;

 always  @(posedge PCLK)
	Ng2360<=Ng2359;

 always  @(posedge PCLK)
	Ng2361<=Ng11575;

 always  @(posedge PCLK)
	Ng2362<=Ng2361;

 always  @(posedge PCLK)
	Ng2363<=Ng11576;

 always  @(posedge PCLK)
	Ng2364<=Ng2363;

 always  @(posedge PCLK)
	Ng2365<=Ng13455;

 always  @(posedge PCLK)
	Ng2366<=Ng2365;

 always  @(posedge PCLK)
	Ng2374<=Ng19048;

 always  @(posedge PCLK)
	Ng2380<=Ng30314;

 always  @(posedge PCLK)
	Ng2373<=Ng27229;

 always  @(posedge PCLK)
	Ng2417<=Ng11578;

 always  @(posedge PCLK)
	Ng2424<=Ng2417;

 always  @(posedge PCLK)
	Ng2425<=Ng11579;

 always  @(posedge PCLK)
	Ng2426<=Ng2425;

 always  @(posedge PCLK)
	Ng2427<=Ng11580;

 always  @(posedge PCLK)
	Ng2428<=Ng2427;

 always  @(posedge PCLK)
	Ng2432<=Ng11581;

 always  @(posedge PCLK)
	Ng2439<=Ng2432;

 always  @(posedge PCLK)
	Ng2440<=Ng11582;

 always  @(posedge PCLK)
	Ng2441<=Ng2440;

 always  @(posedge PCLK)
	Ng2442<=Ng11583;

 always  @(posedge PCLK)
	Ng2443<=Ng2442;

 always  @(posedge PCLK)
	Ng2447<=Ng11584;

 always  @(posedge PCLK)
	Ng2454<=Ng2447;

 always  @(posedge PCLK)
	Ng2455<=Ng11585;

 always  @(posedge PCLK)
	Ng2456<=Ng2455;

 always  @(posedge PCLK)
	Ng2457<=Ng11586;

 always  @(posedge PCLK)
	Ng2458<=Ng2457;

 always  @(posedge PCLK)
	Ng2462<=Ng11587;

 always  @(posedge PCLK)
	Ng2469<=Ng2462;

 always  @(posedge PCLK)
	Ng2470<=Ng11588;

 always  @(posedge PCLK)
	Ng2471<=Ng2470;

 always  @(posedge PCLK)
	Ng2472<=Ng11589;

 always  @(posedge PCLK)
	Ng2399<=Ng2472;

 always  @(posedge PCLK)
	Ng2628<=Ng23274;

 always  @(posedge PCLK)
	Ng2631<=Ng20568;

 always  @(posedge PCLK)
	Ng2584<=Ng20569;

 always  @(posedge PCLK)
	Ng2587<=Ng16473;

 always  @(posedge PCLK)
	Ng2597<=Ng2587;

 always  @(posedge PCLK)
	Ng2598<=Ng2597;

 always  @(posedge PCLK)
	Ng2638<=Ng11593;

 always  @(posedge PCLK)
	Ng2643<=Ng2638;

 always  @(posedge PCLK)
	Ng2644<=Ng11596;

 always  @(posedge PCLK)
	Ng2645<=Ng2644;

 always  @(posedge PCLK)
	Ng2646<=Ng11597;

 always  @(posedge PCLK)
	Ng2647<=Ng2646;

 always  @(posedge PCLK)
	Ng2648<=Ng11598;

 always  @(posedge PCLK)
	Ng2639<=Ng2648;

 always  @(posedge PCLK)
	Ng2640<=Ng11594;

 always  @(posedge PCLK)
	Ng2641<=Ng2640;

 always  @(posedge PCLK)
	Ng2642<=Ng11595;

 always  @(posedge PCLK)
	Ng2564<=Ng2642;

 always  @(posedge PCLK)
	Ng2561<=Ng24415;

 always  @(posedge PCLK)
	Ng2562<=Ng24416;

 always  @(posedge PCLK)
	Ng2563<=Ng24417;

 always  @(posedge PCLK)
	Ng11593<=Ng25172;

 always  @(posedge PCLK)
	Ng11596<=Ng25164;

 always  @(posedge PCLK)
	Ng11597<=Ng25165;

 always  @(posedge PCLK)
	Ng2552<=Ng25169;

 always  @(posedge PCLK)
	Ng2553<=Ng25170;

 always  @(posedge PCLK)
	Ng2554<=Ng25171;

 always  @(posedge PCLK)
	Ng2555<=Ng24412;

 always  @(posedge PCLK)
	Ng2559<=Ng24413;

 always  @(posedge PCLK)
	Ng2539<=Ng24414;

 always  @(posedge PCLK)
	Ng11598<=Ng25166;

 always  @(posedge PCLK)
	Ng11594<=Ng25167;

 always  @(posedge PCLK)
	Ng11595<=Ng25168;

 always  @(posedge PCLK)
	Ng2602<=Ng16474;

 always  @(posedge PCLK)
	Ng2609<=Ng2602;

 always  @(posedge PCLK)
	Ng2616<=Ng2609;

 always  @(posedge PCLK)
	Ng2617<=Ng19057;

 always  @(posedge PCLK)
	Ng2618<=Ng2617;

 always  @(posedge PCLK)
	Ng2622<=Ng30325;

 always  @(posedge PCLK)
	Ng2623<=Ng19058;

 always  @(posedge PCLK)
	Ng8311<=Ng2623;

 always  @(posedge PCLK)
	Ng2632<=Ng19059;

 always  @(posedge PCLK)
	Ng2633<=Ng2632;

 always  @(posedge PCLK)
	Ng2650<=Ng28297;

 always  @(posedge PCLK)
	Ng2651<=Ng28298;

 always  @(posedge PCLK)
	Ng2649<=Ng28299;

 always  @(posedge PCLK)
	Ng2653<=Ng28300;

 always  @(posedge PCLK)
	Ng2654<=Ng28301;

 always  @(posedge PCLK)
	Ng2652<=Ng28302;

 always  @(posedge PCLK)
	Ng2656<=Ng28303;

 always  @(posedge PCLK)
	Ng2657<=Ng28304;

 always  @(posedge PCLK)
	Ng2655<=Ng28305;

 always  @(posedge PCLK)
	Ng2659<=Ng28306;

 always  @(posedge PCLK)
	Ng2660<=Ng28307;

 always  @(posedge PCLK)
	Ng2658<=Ng28308;

 always  @(posedge PCLK)
	Ng2661<=Ng26012;

 always  @(posedge PCLK)
	Ng2664<=Ng26013;

 always  @(posedge PCLK)
	Ng2667<=Ng26014;

 always  @(posedge PCLK)
	Ng2670<=Ng26015;

 always  @(posedge PCLK)
	Ng2673<=Ng26016;

 always  @(posedge PCLK)
	Ng2676<=Ng26017;

 always  @(posedge PCLK)
	Ng2688<=Ng29159;

 always  @(posedge PCLK)
	Ng2691<=Ng29160;

 always  @(posedge PCLK)
	Ng2694<=Ng29161;

 always  @(posedge PCLK)
	Ng2679<=Ng29156;

 always  @(posedge PCLK)
	Ng2682<=Ng29157;

 always  @(posedge PCLK)
	Ng2685<=Ng29158;

 always  @(posedge PCLK)
	Ng2565<=Ng27233;

 always  @(posedge PCLK)
	Ng2568<=Ng27234;

 always  @(posedge PCLK)
	Ng2571<=Ng27235;

 always  @(posedge PCLK)
	Ng2580<=Ng8311;

 always  @(posedge PCLK)
	Ng2581<=Ng24418;

 always  @(posedge PCLK)
	Pg16437<=Ng30320;

 always  @(posedge PCLK)
	Ng2599<=Pg16437;

 always  @(posedge PCLK)
	Ng2603<=Ng13458;

 always  @(posedge PCLK)
	Ng2604<=Ng13459;

 always  @(posedge PCLK)
	Ng2605<=Ng13460;

 always  @(posedge PCLK)
	Ng2606<=Ng13461;

 always  @(posedge PCLK)
	Ng2607<=Ng13462;

 always  @(posedge PCLK)
	Ng2608<=Ng13463;

 always  @(posedge PCLK)
	Ng2610<=Ng13464;

 always  @(posedge PCLK)
	Ng2611<=Ng13465;

 always  @(posedge PCLK)
	Ng2612<=Ng26011;

 always  @(posedge PCLK)
	Ng2615<=Ng13466;

 always  @(posedge PCLK)
	Ng2704<=Ng20570;

 always  @(posedge PCLK)
	Ng2733<=Ng21946;

 always  @(posedge PCLK)
	Ng2714<=Ng23275;

 always  @(posedge PCLK)
	Ng2707<=Ng24419;

 always  @(posedge PCLK)
	Ng2727<=Ng25173;

 always  @(posedge PCLK)
	Ng2720<=Ng26018;

 always  @(posedge PCLK)
	Ng2734<=Ng26742;

 always  @(posedge PCLK)
	Ng2746<=Ng27236;

 always  @(posedge PCLK)
	Ng2740<=Ng27714;

 always  @(posedge PCLK)
	Ng2753<=Ng28309;

 always  @(posedge PCLK)
	Ng2760<=Ng28692;

 always  @(posedge PCLK)
	Ng2766<=Ng29162;

 always  @(posedge PCLK)
	Ng2773<=Ng23276;

 always  @(posedge PCLK)
	Ng2774<=Ng23277;

 always  @(posedge PCLK)
	Ng2772<=Ng23278;

 always  @(posedge PCLK)
	Ng2776<=Ng23279;

 always  @(posedge PCLK)
	Ng2777<=Ng23280;

 always  @(posedge PCLK)
	Ng2775<=Ng23281;

 always  @(posedge PCLK)
	Ng2779<=Ng23282;

 always  @(posedge PCLK)
	Ng2780<=Ng23283;

 always  @(posedge PCLK)
	Ng2778<=Ng23284;

 always  @(posedge PCLK)
	Ng2782<=Ng23285;

 always  @(posedge PCLK)
	Ng2783<=Ng23286;

 always  @(posedge PCLK)
	Ng2781<=Ng23287;

 always  @(posedge PCLK)
	Ng2785<=Ng23288;

 always  @(posedge PCLK)
	Ng2786<=Ng23289;

 always  @(posedge PCLK)
	Ng2784<=Ng23290;

 always  @(posedge PCLK)
	Ng2788<=Ng23291;

 always  @(posedge PCLK)
	Ng2789<=Ng23292;

 always  @(posedge PCLK)
	Ng2787<=Ng23293;

 always  @(posedge PCLK)
	Ng2791<=Ng23294;

 always  @(posedge PCLK)
	Ng2792<=Ng23295;

 always  @(posedge PCLK)
	Ng2790<=Ng23296;

 always  @(posedge PCLK)
	Ng2794<=Ng23297;

 always  @(posedge PCLK)
	Ng2795<=Ng23298;

 always  @(posedge PCLK)
	Ng2793<=Ng23299;

 always  @(posedge PCLK)
	Ng2797<=Ng23300;

 always  @(posedge PCLK)
	Ng2798<=Ng23301;

 always  @(posedge PCLK)
	Ng2796<=Ng23302;

 always  @(posedge PCLK)
	Ng2800<=Ng23303;

 always  @(posedge PCLK)
	Ng2801<=Ng23304;

 always  @(posedge PCLK)
	Ng2799<=Ng23305;

 always  @(posedge PCLK)
	Ng2803<=Ng23306;

 always  @(posedge PCLK)
	Ng2804<=Ng23307;

 always  @(posedge PCLK)
	Ng2802<=Ng23308;

 always  @(posedge PCLK)
	Ng2806<=Ng23309;

 always  @(posedge PCLK)
	Ng2807<=Ng23310;

 always  @(posedge PCLK)
	Ng2805<=Ng23311;

 always  @(posedge PCLK)
	Ng2809<=Ng26743;

 always  @(posedge PCLK)
	Ng2810<=Ng26744;

 always  @(posedge PCLK)
	Ng2808<=Ng26745;

 always  @(posedge PCLK)
	Ng2812<=Ng24420;

 always  @(posedge PCLK)
	Ng2813<=Ng24421;

 always  @(posedge PCLK)
	Ng2811<=Ng24422;

 always  @(posedge PCLK)
	Ng3054<=Ng23317;

 always  @(posedge PCLK)
	Ng3079<=Ng23318;

 always  @(posedge PCLK)
	Ng13475<=Ng21965;

 always  @(posedge PCLK)
	Ng3043<=Ng29453;

 always  @(posedge PCLK)
	Ng3044<=Ng29454;

 always  @(posedge PCLK)
	Ng3045<=Ng29455;

 always  @(posedge PCLK)
	Ng3046<=Ng29456;

 always  @(posedge PCLK)
	Ng3047<=Ng29457;

 always  @(posedge PCLK)
	Ng3048<=Ng29458;

 always  @(posedge PCLK)
	Ng3049<=Ng29459;

 always  @(posedge PCLK)
	Ng3050<=Ng29460;

 always  @(posedge PCLK)
	Ng3051<=Ng29655;

 always  @(posedge PCLK)
	Ng3052<=Ng29972;

 always  @(posedge PCLK)
	Ng3053<=Ng29973;

 always  @(posedge PCLK)
	Ng3055<=Ng29974;

 always  @(posedge PCLK)
	Ng3056<=Ng29975;

 always  @(posedge PCLK)
	Ng3057<=Ng29976;

 always  @(posedge PCLK)
	Ng3058<=Ng29977;

 always  @(posedge PCLK)
	Ng3059<=Ng29978;

 always  @(posedge PCLK)
	Ng3060<=Ng29979;

 always  @(posedge PCLK)
	Ng3061<=Ng30119;

 always  @(posedge PCLK)
	Ng3062<=Ng30908;

 always  @(posedge PCLK)
	Ng3063<=Ng30909;

 always  @(posedge PCLK)
	Ng3064<=Ng30910;

 always  @(posedge PCLK)
	Ng3065<=Ng30911;

 always  @(posedge PCLK)
	Ng3066<=Ng30912;

 always  @(posedge PCLK)
	Ng3067<=Ng30913;

 always  @(posedge PCLK)
	Ng3068<=Ng30914;

 always  @(posedge PCLK)
	Ng3069<=Ng30915;

 always  @(posedge PCLK)
	Ng3070<=Ng30940;

 always  @(posedge PCLK)
	Ng3071<=Ng30980;

 always  @(posedge PCLK)
	Ng3072<=Ng30981;

 always  @(posedge PCLK)
	Ng3073<=Ng30982;

 always  @(posedge PCLK)
	Ng3074<=Ng30983;

 always  @(posedge PCLK)
	Ng3075<=Ng30984;

 always  @(posedge PCLK)
	Ng3076<=Ng30985;

 always  @(posedge PCLK)
	Ng3077<=Ng30986;

 always  @(posedge PCLK)
	Ng3078<=Ng30987;

 always  @(posedge PCLK)
	Ng2997<=Ng30989;

 always  @(posedge PCLK)
	Ng2993<=Ng26748;

 always  @(posedge PCLK)
	Ng2998<=Ng27238;

 always  @(posedge PCLK)
	Ng3006<=Ng25177;

 always  @(posedge PCLK)
	Ng3002<=Ng26021;

 always  @(posedge PCLK)
	Ng3013<=Ng26750;

 always  @(posedge PCLK)
	Ng3010<=Ng27239;

 always  @(posedge PCLK)
	Ng3024<=Ng27716;

 always  @(posedge PCLK)
	Ng3018<=Ng24425;

 always  @(posedge PCLK)
	Ng3028<=Ng25176;

 always  @(posedge PCLK)
	Ng3036<=Ng26022;

 always  @(posedge PCLK)
	Ng3032<=Ng26749;

 always  @(posedge PCLK)
	Pg5388<=Pg3234;

 always  @(posedge PCLK)
	Ng2986<=Pg5388;

 always  @(posedge PCLK)
	Ng2987<=Pg16496;

 always  @(posedge PCLK)
	Pg8275<=Ng20595;

 always  @(posedge PCLK)
	Pg8274<=Ng20596;

 always  @(posedge PCLK)
	Pg8273<=Ng20597;

 always  @(posedge PCLK)
	Pg8272<=Ng20598;

 always  @(posedge PCLK)
	Pg8268<=Ng20599;

 always  @(posedge PCLK)
	Pg8269<=Ng20600;

 always  @(posedge PCLK)
	Pg8270<=Ng20601;

 always  @(posedge PCLK)
	Pg8271<=Ng20602;

 always  @(posedge PCLK)
	Ng3083<=Ng20603;

 always  @(posedge PCLK)
	Pg8267<=Ng20604;

 always  @(posedge PCLK)
	Ng2992<=Ng21966;

 always  @(posedge PCLK)
	Pg8266<=Ng20605;

 always  @(posedge PCLK)
	Pg8265<=Ng20606;

 always  @(posedge PCLK)
	Pg8264<=Ng20607;

 always  @(posedge PCLK)
	Pg8262<=Ng20608;

 always  @(posedge PCLK)
	Pg8263<=Ng20589;

 always  @(posedge PCLK)
	Pg8260<=Ng20590;

 always  @(posedge PCLK)
	Pg8261<=Ng20591;

 always  @(posedge PCLK)
	Pg8259<=Ng20592;

 always  @(posedge PCLK)
	Ng2990<=Ng20593;

 always  @(posedge PCLK)
	Ng2991<=Ng21964;

 always  @(posedge PCLK)
	Pg8258<=Ng20594;

 assign Pg27380 = ( (~ Ng29656) ) ;
 assign Pg26149 = ( (~ n1770) ) ;
 assign Pg26135 = ( (~ Ng29166) ) ;
 assign Pg26104 = ( (~ n1778) ) ;
 assign Pg25489 = ( (~ n3323) ) ;
 assign wire1521 = ( (~ Pg3233) ) | ( Pg3230 ) ;
 assign Pg25435 = ( (~ Ng28696) ) ;
 assign Pg24734 = ( (~ Ng28313) ) ;
 assign Pg16496 = ( (~ n188) ) ;
 assign n1139 = ( (~ Pg8269)  &  Pg8268 ) | ( Pg8269  &  (~ Pg8268) ) ;
 assign n1138 = ( (~ Pg8271)  &  Pg8270 ) | ( Pg8271  &  (~ Pg8270) ) ;
 assign n1137 = ( (~ n1139)  &  n1138 ) | ( n1139  &  (~ n1138) ) ;
 assign n1142 = ( (~ Pg8262)  &  Pg8264 ) | ( Pg8262  &  (~ Pg8264) ) ;
 assign n1141 = ( (~ Pg8265)  &  Pg8266 ) | ( Pg8265  &  (~ Pg8266) ) ;
 assign n1140 = ( (~ n1142)  &  n1141 ) | ( n1142  &  (~ n1141) ) ;
 assign n1145 = ( (~ Pg8259)  &  Pg8261 ) | ( Pg8259  &  (~ Pg8261) ) ;
 assign n1144 = ( (~ Pg8260)  &  Pg8263 ) | ( Pg8260  &  (~ Pg8263) ) ;
 assign n1143 = ( (~ n1145)  &  n1144 ) | ( n1145  &  (~ n1144) ) ;
 assign n1148 = ( (~ Pg8272)  &  Pg8273 ) | ( Pg8272  &  (~ Pg8273) ) ;
 assign n1147 = ( (~ Pg8275)  &  Pg8274 ) | ( Pg8275  &  (~ Pg8274) ) ;
 assign n1146 = ( (~ n1148)  &  n1147 ) | ( n1148  &  (~ n1147) ) ;
 assign n69 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng324) ) | ( (~ Ng1315)  &  (~ Ng394) ) | ( (~ Ng324)  &  (~ Ng394) ) ;
 assign n66 = ( (~ wire1603)  &  n69 ) | ( n69  &  (~ Ng396) ) ;
 assign n72 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng383) ) | ( (~ Ng1315)  &  (~ Ng379) ) | ( (~ Ng383)  &  (~ Ng379) ) ;
 assign n70 = ( (~ wire1603)  &  n72 ) | ( n72  &  (~ Ng381) ) ;
 assign n75 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1011) ) | ( (~ Ng1315)  &  (~ Ng1081) ) | ( (~ Ng1011)  &  (~ Ng1081) ) ;
 assign n73 = ( (~ wire1603)  &  n75 ) | ( n75  &  (~ Ng1083) ) ;
 assign n78 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng368) ) | ( (~ Ng1315)  &  (~ Ng364) ) | ( (~ Ng368)  &  (~ Ng364) ) ;
 assign n76 = ( (~ wire1603)  &  n78 ) | ( n78  &  (~ Ng366) ) ;
 assign n81 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1070) ) | ( (~ Ng1315)  &  (~ Ng1066) ) | ( (~ Ng1070)  &  (~ Ng1066) ) ;
 assign n79 = ( (~ wire1603)  &  n81 ) | ( n81  &  (~ Ng1068) ) ;
 assign n84 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1705) ) | ( (~ Ng1315)  &  (~ Ng1775) ) | ( (~ Ng1705)  &  (~ Ng1775) ) ;
 assign n82 = ( (~ wire1603)  &  n84 ) | ( n84  &  (~ Ng1777) ) ;
 assign n87 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng353) ) | ( (~ Ng1315)  &  (~ Ng349) ) | ( (~ Ng353)  &  (~ Ng349) ) ;
 assign n85 = ( (~ wire1603)  &  n87 ) | ( n87  &  (~ Ng351) ) ;
 assign n90 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1055) ) | ( (~ Ng1315)  &  (~ Ng1051) ) | ( (~ Ng1055)  &  (~ Ng1051) ) ;
 assign n88 = ( (~ wire1603)  &  n90 ) | ( n90  &  (~ Ng1053) ) ;
 assign n93 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1764) ) | ( (~ Ng1315)  &  (~ Ng1760) ) | ( (~ Ng1764)  &  (~ Ng1760) ) ;
 assign n91 = ( (~ wire1603)  &  n93 ) | ( n93  &  (~ Ng1762) ) ;
 assign n96 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2399) ) | ( (~ Ng1315)  &  (~ Ng2469) ) | ( (~ Ng2399)  &  (~ Ng2469) ) ;
 assign n94 = ( (~ wire1603)  &  n96 ) | ( n96  &  (~ Ng2471) ) ;
 assign n99 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1040) ) | ( (~ Ng1315)  &  (~ Ng1036) ) | ( (~ Ng1040)  &  (~ Ng1036) ) ;
 assign n97 = ( (~ wire1603)  &  n99 ) | ( n99  &  (~ Ng1038) ) ;
 assign n102 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1749) ) | ( (~ Ng1315)  &  (~ Ng1745) ) | ( (~ Ng1749)  &  (~ Ng1745) ) ;
 assign n100 = ( (~ wire1603)  &  n102 ) | ( n102  &  (~ Ng1747) ) ;
 assign n105 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2458) ) | ( (~ Ng1315)  &  (~ Ng2454) ) | ( (~ Ng2458)  &  (~ Ng2454) ) ;
 assign n103 = ( (~ wire1603)  &  n105 ) | ( n105  &  (~ Ng2456) ) ;
 assign n108 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1734) ) | ( (~ Ng1315)  &  (~ Ng1730) ) | ( (~ Ng1734)  &  (~ Ng1730) ) ;
 assign n106 = ( (~ wire1603)  &  n108 ) | ( n108  &  (~ Ng1732) ) ;
 assign n111 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2443) ) | ( (~ Ng1315)  &  (~ Ng2439) ) | ( (~ Ng2443)  &  (~ Ng2439) ) ;
 assign n109 = ( (~ wire1603)  &  n111 ) | ( n111  &  (~ Ng2441) ) ;
 assign n114 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2428) ) | ( (~ Ng1315)  &  (~ Ng2424) ) | ( (~ Ng2428)  &  (~ Ng2424) ) ;
 assign n112 = ( (~ wire1603)  &  n114 ) | ( n114  &  (~ Ng2426) ) ;
 assign n117 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng496) ) | ( (~ Ng1315)  &  (~ Ng490) ) | ( (~ Ng496)  &  (~ Ng490) ) ;
 assign n115 = ( (~ wire1603)  &  n117 ) | ( n117  &  (~ Ng493) ) ;
 assign n120 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1183) ) | ( (~ Ng1315)  &  (~ Ng1177) ) | ( (~ Ng1183)  &  (~ Ng1177) ) ;
 assign n118 = ( (~ wire1603)  &  n120 ) | ( n120  &  (~ Ng1180) ) ;
 assign n123 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1877) ) | ( (~ Ng1315)  &  (~ Ng1871) ) | ( (~ Ng1877)  &  (~ Ng1871) ) ;
 assign n121 = ( (~ wire1603)  &  n123 ) | ( n123  &  (~ Ng1874) ) ;
 assign n126 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2571) ) | ( (~ Ng1315)  &  (~ Ng2565) ) | ( (~ Ng2571)  &  (~ Ng2565) ) ;
 assign n124 = ( (~ wire1603)  &  n126 ) | ( n126  &  (~ Ng2568) ) ;
 assign n129 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ Ng853)  &  Ng448 ) | ( (~ wire1612)  &  Ng447 ) | ( Ng448  &  Ng447 ) ;
 assign n127 = ( (~ wire1594)  &  n129 ) | ( n129  &  Ng449 ) ;
 assign n131 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng402 ) | ( (~ Ng853)  &  Ng403 ) | ( Ng402  &  Ng403 ) ;
 assign n130 = ( (~ wire1594)  &  n131 ) | ( n131  &  Ng404 ) ;
 assign n133 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng479 ) | ( (~ wire1605)  &  Ng477 ) | ( Ng479  &  Ng477 ) ;
 assign Ng19021 = ( (~ Ng1315)  &  n133 ) | ( n133  &  Ng478 ) ;
 assign n134 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng464 ) | ( (~ wire1605)  &  Ng480 ) | ( Ng464  &  Ng480 ) ;
 assign Ng19022 = ( (~ Ng1315)  &  n134 ) | ( n134  &  Ng484 ) ;
 assign n136 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ Ng853)  &  Ng1135 ) | ( (~ wire1612)  &  Ng1134 ) | ( Ng1135  &  Ng1134 ) ;
 assign n135 = ( (~ wire1594)  &  n136 ) | ( n136  &  Ng1136 ) ;
 assign n138 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1089 ) | ( (~ Ng853)  &  Ng1090 ) | ( Ng1089  &  Ng1090 ) ;
 assign n137 = ( (~ wire1594)  &  n138 ) | ( n138  &  Ng1091 ) ;
 assign n139 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng1166 ) | ( (~ wire1605)  &  Ng1164 ) | ( Ng1166  &  Ng1164 ) ;
 assign Ng19033 = ( (~ Ng1315)  &  n139 ) | ( n139  &  Ng1165 ) ;
 assign n140 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng488 ) | ( (~ wire1605)  &  Ng486 ) | ( Ng488  &  Ng486 ) ;
 assign Ng19023 = ( (~ Ng1315)  &  n140 ) | ( n140  &  Ng487 ) ;
 assign n141 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng1151 ) | ( (~ wire1605)  &  Ng1167 ) | ( Ng1151  &  Ng1167 ) ;
 assign Ng19034 = ( (~ Ng1315)  &  n141 ) | ( n141  &  Ng1171 ) ;
 assign n143 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ Ng853)  &  Ng1829 ) | ( (~ wire1612)  &  Ng1828 ) | ( Ng1829  &  Ng1828 ) ;
 assign n142 = ( (~ wire1594)  &  n143 ) | ( n143  &  Ng1830 ) ;
 assign n145 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1783 ) | ( (~ Ng853)  &  Ng1784 ) | ( Ng1783  &  Ng1784 ) ;
 assign n144 = ( (~ wire1594)  &  n145 ) | ( n145  &  Ng1785 ) ;
 assign n146 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng1860 ) | ( (~ wire1605)  &  Ng1858 ) | ( Ng1860  &  Ng1858 ) ;
 assign Ng19045 = ( (~ Ng1315)  &  n146 ) | ( n146  &  Ng1859 ) ;
 assign n148 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng573) ) | ( (~ Ng1315)  &  (~ Ng569) ) | ( (~ Ng573)  &  (~ Ng569) ) ;
 assign Ng16467 = ( (~ wire1603)  &  n148 ) | ( n148  &  (~ Ng571) ) ;
 assign n149 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng1175 ) | ( (~ wire1605)  &  Ng1173 ) | ( Ng1175  &  Ng1173 ) ;
 assign Ng19035 = ( (~ Ng1315)  &  n149 ) | ( n149  &  Ng1174 ) ;
 assign n150 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng1845 ) | ( (~ wire1605)  &  Ng1861 ) | ( Ng1845  &  Ng1861 ) ;
 assign Ng19046 = ( (~ Ng1315)  &  n150 ) | ( n150  &  Ng1865 ) ;
 assign n152 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ Ng853)  &  Ng2523 ) | ( (~ wire1612)  &  Ng2522 ) | ( Ng2523  &  Ng2522 ) ;
 assign n151 = ( (~ wire1594)  &  n152 ) | ( n152  &  Ng2524 ) ;
 assign n154 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2477 ) | ( (~ Ng853)  &  Ng2478 ) | ( Ng2477  &  Ng2478 ) ;
 assign n153 = ( (~ wire1594)  &  n154 ) | ( n154  &  Ng2479 ) ;
 assign n155 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng2554 ) | ( (~ wire1605)  &  Ng2552 ) | ( Ng2554  &  Ng2552 ) ;
 assign Ng19057 = ( (~ Ng1315)  &  n155 ) | ( n155  &  Ng2553 ) ;
 assign n157 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1259) ) | ( (~ Ng1315)  &  (~ Ng1255) ) | ( (~ Ng1259)  &  (~ Ng1255) ) ;
 assign Ng16469 = ( (~ wire1603)  &  n157 ) | ( n157  &  (~ Ng1257) ) ;
 assign n158 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng1869 ) | ( (~ wire1605)  &  Ng1867 ) | ( Ng1869  &  Ng1867 ) ;
 assign Ng19047 = ( (~ Ng1315)  &  n158 ) | ( n158  &  Ng1868 ) ;
 assign n159 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng2539 ) | ( (~ wire1605)  &  Ng2555 ) | ( Ng2539  &  Ng2555 ) ;
 assign Ng19058 = ( (~ Ng1315)  &  n159 ) | ( n159  &  Ng2559 ) ;
 assign n161 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng321 ) | ( (~ Ng853)  &  Ng322 ) | ( Ng321  &  Ng322 ) ;
 assign n160 = ( (~ wire1594)  &  n161 ) | ( n161  &  Ng323 ) ;
 assign n163 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1953) ) | ( (~ Ng1315)  &  (~ Ng1949) ) | ( (~ Ng1953)  &  (~ Ng1949) ) ;
 assign Ng16471 = ( (~ wire1603)  &  n163 ) | ( n163  &  (~ Ng1951) ) ;
 assign n164 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1603)  &  Ng2563 ) | ( (~ wire1605)  &  Ng2561 ) | ( Ng2563  &  Ng2561 ) ;
 assign Ng19059 = ( (~ Ng1315)  &  n164 ) | ( n164  &  Ng2562 ) ;
 assign n166 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng489) ) | ( (~ Ng1315)  &  (~ Ng565) ) | ( (~ Ng489)  &  (~ Ng565) ) ;
 assign Ng16468 = ( (~ wire1603)  &  n166 ) | ( n166  &  (~ Ng567) ) ;
 assign n168 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1008 ) | ( (~ Ng853)  &  Ng1009 ) | ( Ng1008  &  Ng1009 ) ;
 assign n167 = ( (~ wire1594)  &  n168 ) | ( n168  &  Ng1010 ) ;
 assign n170 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2647) ) | ( (~ Ng1315)  &  (~ Ng2643) ) | ( (~ Ng2647)  &  (~ Ng2643) ) ;
 assign Ng16473 = ( (~ wire1603)  &  n170 ) | ( n170  &  (~ Ng2645) ) ;
 assign n172 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1176) ) | ( (~ Ng1315)  &  (~ Ng1251) ) | ( (~ Ng1176)  &  (~ Ng1251) ) ;
 assign Ng16470 = ( (~ wire1603)  &  n172 ) | ( n172  &  (~ Ng1253) ) ;
 assign n174 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1702 ) | ( (~ Ng853)  &  Ng1703 ) | ( Ng1702  &  Ng1703 ) ;
 assign n173 = ( (~ wire1594)  &  n174 ) | ( n174  &  Ng1704 ) ;
 assign n176 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1870) ) | ( (~ Ng1315)  &  (~ Ng1945) ) | ( (~ Ng1870)  &  (~ Ng1945) ) ;
 assign Ng16472 = ( (~ wire1603)  &  n176 ) | ( n176  &  (~ Ng1947) ) ;
 assign n178 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2396 ) | ( (~ Ng853)  &  Ng2397 ) | ( Ng2396  &  Ng2397 ) ;
 assign n177 = ( (~ wire1594)  &  n178 ) | ( n178  &  Ng2398 ) ;
 assign n180 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2564) ) | ( (~ Ng1315)  &  (~ Ng2639) ) | ( (~ Ng2564)  &  (~ Ng2639) ) ;
 assign Ng16474 = ( (~ wire1603)  &  n180 ) | ( n180  &  (~ Ng2641) ) ;
 assign n183 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng141 ) | ( (~ Ng853)  &  Ng143 ) | ( Ng141  &  Ng143 ) ;
 assign n181 = ( (~ wire1612)  &  n183 ) | ( n183  &  Ng142 ) ;
 assign n185 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng144 ) | ( (~ Ng853)  &  Ng146 ) | ( Ng144  &  Ng146 ) ;
 assign n184 = ( (~ wire1612)  &  n185 ) | ( n185  &  Ng145 ) ;
 assign n187 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng829 ) | ( (~ Ng853)  &  Ng831 ) | ( Ng829  &  Ng831 ) ;
 assign n186 = ( (~ wire1612)  &  n187 ) | ( n187  &  Ng830 ) ;
 assign n188 = ( (~ Pg5388)  &  Ng2987 ) | ( Ng2987  &  Ng2986 ) ;
 assign n190 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng147 ) | ( (~ Ng853)  &  Ng149 ) | ( Ng147  &  Ng149 ) ;
 assign n189 = ( (~ wire1612)  &  n190 ) | ( n190  &  Ng148 ) ;
 assign n192 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng832 ) | ( (~ Ng853)  &  Ng834 ) | ( Ng832  &  Ng834 ) ;
 assign n191 = ( (~ wire1612)  &  n192 ) | ( n192  &  Ng833 ) ;
 assign n194 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng1523 ) | ( (~ Ng853)  &  Ng1525 ) | ( Ng1523  &  Ng1525 ) ;
 assign n193 = ( (~ wire1612)  &  n194 ) | ( n194  &  Ng1524 ) ;
 assign n196 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng150 ) | ( (~ Ng853)  &  Ng152 ) | ( Ng150  &  Ng152 ) ;
 assign n195 = ( (~ wire1612)  &  n196 ) | ( n196  &  Ng151 ) ;
 assign n199 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ Ng853)  &  (~ Ng216) ) | ( (~ wire1594)  &  (~ Ng219) ) | ( (~ Ng216)  &  (~ Ng219) ) ;
 assign n197 = ( (~ wire1612)  &  n199 ) | ( n199  &  (~ Ng213) ) ;
 assign n201 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng835 ) | ( (~ Ng853)  &  Ng837 ) | ( Ng835  &  Ng837 ) ;
 assign n200 = ( (~ wire1612)  &  n201 ) | ( n201  &  Ng836 ) ;
 assign n203 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng1526 ) | ( (~ Ng853)  &  Ng1528 ) | ( Ng1526  &  Ng1528 ) ;
 assign n202 = ( (~ wire1612)  &  n203 ) | ( n203  &  Ng1527 ) ;
 assign n205 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng2217 ) | ( (~ Ng853)  &  Ng2219 ) | ( Ng2217  &  Ng2219 ) ;
 assign n204 = ( (~ wire1612)  &  n205 ) | ( n205  &  Ng2218 ) ;
 assign n207 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng153 ) | ( (~ Ng853)  &  Ng154 ) | ( Ng153  &  Ng154 ) ;
 assign n206 = ( (~ wire1594)  &  n207 ) | ( n207  &  Ng155 ) ;
 assign n211 = ( (~ wire1594)  &  (~ wire1612) ) | ( (~ wire1594)  &  (~ Ng222) ) | ( (~ wire1612)  &  (~ Ng225) ) | ( (~ Ng222)  &  (~ Ng225) ) ;
 assign n208 = ( (~ Ng853)  &  n211 ) | ( n211  &  (~ Ng228) ) ;
 assign n213 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng838 ) | ( (~ Ng853)  &  Ng839 ) | ( Ng838  &  Ng839 ) ;
 assign n212 = ( (~ wire1594)  &  n213 ) | ( n213  &  Ng840 ) ;
 assign n216 = ( (~ wire1594)  &  (~ wire1612) ) | ( (~ wire1594)  &  (~ Ng900) ) | ( (~ wire1612)  &  (~ Ng903) ) | ( (~ Ng900)  &  (~ Ng903) ) ;
 assign n214 = ( (~ Ng853)  &  n216 ) | ( n216  &  (~ Ng906) ) ;
 assign n218 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1529 ) | ( (~ Ng853)  &  Ng1530 ) | ( Ng1529  &  Ng1530 ) ;
 assign n217 = ( (~ wire1594)  &  n218 ) | ( n218  &  Ng1531 ) ;
 assign n220 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2220 ) | ( (~ Ng853)  &  Ng2221 ) | ( Ng2220  &  Ng2221 ) ;
 assign n219 = ( (~ wire1594)  &  n220 ) | ( n220  &  Ng2222 ) ;
 assign n222 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng156 ) | ( (~ Ng853)  &  Ng157 ) | ( Ng156  &  Ng157 ) ;
 assign n221 = ( (~ wire1594)  &  n222 ) | ( n222  &  Ng158 ) ;
 assign n225 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng237) ) | ( (~ Ng853)  &  (~ Ng231) ) | ( (~ Ng237)  &  (~ Ng231) ) ;
 assign n223 = ( (~ wire1594)  &  n225 ) | ( n225  &  (~ Ng234) ) ;
 assign n227 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng698 ) | ( (~ Ng1315)  &  Ng699 ) | ( Ng698  &  Ng699 ) ;
 assign n226 = ( (~ wire1603)  &  n227 ) | ( n227  &  Ng700 ) ;
 assign n229 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng725 ) | ( (~ Ng1315)  &  Ng726 ) | ( Ng725  &  Ng726 ) ;
 assign n228 = ( (~ wire1603)  &  n229 ) | ( n229  &  Ng727 ) ;
 assign n231 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng841 ) | ( (~ Ng853)  &  Ng842 ) | ( Ng841  &  Ng842 ) ;
 assign n230 = ( (~ wire1594)  &  n231 ) | ( n231  &  Ng843 ) ;
 assign n234 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng915) ) | ( (~ Ng853)  &  (~ Ng909) ) | ( (~ Ng915)  &  (~ Ng909) ) ;
 assign n232 = ( (~ wire1594)  &  n234 ) | ( n234  &  (~ Ng912) ) ;
 assign n236 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1532 ) | ( (~ Ng853)  &  Ng1533 ) | ( Ng1532  &  Ng1533 ) ;
 assign n235 = ( (~ wire1594)  &  n236 ) | ( n236  &  Ng1534 ) ;
 assign n239 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1600) ) | ( (~ Ng853)  &  (~ Ng1594) ) | ( (~ Ng1600)  &  (~ Ng1594) ) ;
 assign n237 = ( (~ wire1594)  &  n239 ) | ( n239  &  (~ Ng1597) ) ;
 assign n241 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2223 ) | ( (~ Ng853)  &  Ng2224 ) | ( Ng2223  &  Ng2224 ) ;
 assign n240 = ( (~ wire1594)  &  n241 ) | ( n241  &  Ng2225 ) ;
 assign n243 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng159 ) | ( (~ Ng853)  &  Ng160 ) | ( Ng159  &  Ng160 ) ;
 assign n242 = ( (~ wire1594)  &  n243 ) | ( n243  &  Ng161 ) ;
 assign n246 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng246) ) | ( (~ Ng853)  &  (~ Ng240) ) | ( (~ Ng246)  &  (~ Ng240) ) ;
 assign n244 = ( (~ wire1594)  &  n246 ) | ( n246  &  (~ Ng243) ) ;
 assign n248 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng701 ) | ( (~ Ng1315)  &  Ng702 ) | ( Ng701  &  Ng702 ) ;
 assign n247 = ( (~ wire1603)  &  n248 ) | ( n248  &  Ng703 ) ;
 assign n250 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng844 ) | ( (~ Ng853)  &  Ng845 ) | ( Ng844  &  Ng845 ) ;
 assign n249 = ( (~ wire1594)  &  n250 ) | ( n250  &  Ng846 ) ;
 assign n253 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng924) ) | ( (~ Ng853)  &  (~ Ng918) ) | ( (~ Ng924)  &  (~ Ng918) ) ;
 assign n251 = ( (~ wire1594)  &  n253 ) | ( n253  &  (~ Ng921) ) ;
 assign n255 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1384 ) | ( (~ Ng1315)  &  Ng1385 ) | ( Ng1384  &  Ng1385 ) ;
 assign n254 = ( (~ wire1603)  &  n255 ) | ( n255  &  Ng1386 ) ;
 assign n257 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1411 ) | ( (~ Ng1315)  &  Ng1412 ) | ( Ng1411  &  Ng1412 ) ;
 assign n256 = ( (~ wire1603)  &  n257 ) | ( n257  &  Ng1413 ) ;
 assign n259 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1535 ) | ( (~ Ng853)  &  Ng1536 ) | ( Ng1535  &  Ng1536 ) ;
 assign n258 = ( (~ wire1594)  &  n259 ) | ( n259  &  Ng1537 ) ;
 assign n262 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1609) ) | ( (~ Ng853)  &  (~ Ng1603) ) | ( (~ Ng1609)  &  (~ Ng1603) ) ;
 assign n260 = ( (~ wire1594)  &  n262 ) | ( n262  &  (~ Ng1606) ) ;
 assign n264 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2226 ) | ( (~ Ng853)  &  Ng2227 ) | ( Ng2226  &  Ng2227 ) ;
 assign n263 = ( (~ wire1594)  &  n264 ) | ( n264  &  Ng2228 ) ;
 assign n267 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2294) ) | ( (~ Ng853)  &  (~ Ng2288) ) | ( (~ Ng2294)  &  (~ Ng2288) ) ;
 assign n265 = ( (~ wire1594)  &  n267 ) | ( n267  &  (~ Ng2291) ) ;
 assign n269 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng129 ) | ( (~ Ng853)  &  Ng130 ) | ( Ng129  &  Ng130 ) ;
 assign n268 = ( (~ wire1594)  &  n269 ) | ( n269  &  Ng131 ) ;
 assign n271 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng162 ) | ( (~ Ng853)  &  Ng163 ) | ( Ng162  &  Ng163 ) ;
 assign n270 = ( (~ wire1594)  &  n271 ) | ( n271  &  Ng164 ) ;
 assign n274 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng255) ) | ( (~ Ng853)  &  (~ Ng249) ) | ( (~ Ng255)  &  (~ Ng249) ) ;
 assign n272 = ( (~ wire1594)  &  n274 ) | ( n274  &  (~ Ng252) ) ;
 assign n276 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng704 ) | ( (~ Ng1315)  &  Ng705 ) | ( Ng704  &  Ng705 ) ;
 assign n275 = ( (~ wire1603)  &  n276 ) | ( n276  &  Ng706 ) ;
 assign n278 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng847 ) | ( (~ Ng853)  &  Ng848 ) | ( Ng847  &  Ng848 ) ;
 assign n277 = ( (~ wire1594)  &  n278 ) | ( n278  &  Ng849 ) ;
 assign n281 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng933) ) | ( (~ Ng853)  &  (~ Ng927) ) | ( (~ Ng933)  &  (~ Ng927) ) ;
 assign n279 = ( (~ wire1594)  &  n281 ) | ( n281  &  (~ Ng930) ) ;
 assign n283 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1387 ) | ( (~ Ng1315)  &  Ng1388 ) | ( Ng1387  &  Ng1388 ) ;
 assign n282 = ( (~ wire1603)  &  n283 ) | ( n283  &  Ng1389 ) ;
 assign n285 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1538 ) | ( (~ Ng853)  &  Ng1539 ) | ( Ng1538  &  Ng1539 ) ;
 assign n284 = ( (~ wire1594)  &  n285 ) | ( n285  &  Ng1540 ) ;
 assign n288 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1618) ) | ( (~ Ng853)  &  (~ Ng1612) ) | ( (~ Ng1618)  &  (~ Ng1612) ) ;
 assign n286 = ( (~ wire1594)  &  n288 ) | ( n288  &  (~ Ng1615) ) ;
 assign n290 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2078 ) | ( (~ Ng1315)  &  Ng2079 ) | ( Ng2078  &  Ng2079 ) ;
 assign n289 = ( (~ wire1603)  &  n290 ) | ( n290  &  Ng2080 ) ;
 assign n292 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2105 ) | ( (~ Ng1315)  &  Ng2106 ) | ( Ng2105  &  Ng2106 ) ;
 assign n291 = ( (~ wire1603)  &  n292 ) | ( n292  &  Ng2107 ) ;
 assign n294 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2229 ) | ( (~ Ng853)  &  Ng2230 ) | ( Ng2229  &  Ng2230 ) ;
 assign n293 = ( (~ wire1594)  &  n294 ) | ( n294  &  Ng2231 ) ;
 assign n297 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2303) ) | ( (~ Ng853)  &  (~ Ng2297) ) | ( (~ Ng2303)  &  (~ Ng2297) ) ;
 assign n295 = ( (~ wire1594)  &  n297 ) | ( n297  &  (~ Ng2300) ) ;
 assign n299 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng132 ) | ( (~ Ng853)  &  Ng133 ) | ( Ng132  &  Ng133 ) ;
 assign n298 = ( (~ wire1594)  &  n299 ) | ( n299  &  Ng134 ) ;
 assign n302 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng264) ) | ( (~ Ng853)  &  (~ Ng258) ) | ( (~ Ng264)  &  (~ Ng258) ) ;
 assign n300 = ( (~ wire1594)  &  n302 ) | ( n302  &  (~ Ng261) ) ;
 assign n304 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11499 ) | ( (~ Ng853)  &  Ng11497 ) | ( Ng11499  &  Ng11497 ) ;
 assign n303 = ( (~ wire1594)  &  n304 ) | ( n304  &  Ng11498 ) ;
 assign n307 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng435) ) | ( (~ Ng853)  &  (~ Ng429) ) | ( (~ Ng435)  &  (~ Ng429) ) ;
 assign n305 = ( (~ wire1594)  &  n307 ) | ( n307  &  (~ Ng432) ) ;
 assign n309 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng707 ) | ( (~ Ng1315)  &  Ng708 ) | ( Ng707  &  Ng708 ) ;
 assign n308 = ( (~ wire1603)  &  n309 ) | ( n309  &  Ng709 ) ;
 assign n311 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng817 ) | ( (~ Ng853)  &  Ng818 ) | ( Ng817  &  Ng818 ) ;
 assign n310 = ( (~ wire1594)  &  n311 ) | ( n311  &  Ng819 ) ;
 assign n313 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng850 ) | ( (~ Ng853)  &  Ng851 ) | ( Ng850  &  Ng851 ) ;
 assign n312 = ( (~ wire1594)  &  n313 ) | ( n313  &  Ng852 ) ;
 assign n316 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng942) ) | ( (~ Ng853)  &  (~ Ng936) ) | ( (~ Ng942)  &  (~ Ng936) ) ;
 assign n314 = ( (~ wire1594)  &  n316 ) | ( n316  &  (~ Ng939) ) ;
 assign n318 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1390 ) | ( (~ Ng1315)  &  Ng1391 ) | ( Ng1390  &  Ng1391 ) ;
 assign n317 = ( (~ wire1603)  &  n318 ) | ( n318  &  Ng1392 ) ;
 assign n320 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1541 ) | ( (~ Ng853)  &  Ng1542 ) | ( Ng1541  &  Ng1542 ) ;
 assign n319 = ( (~ wire1594)  &  n320 ) | ( n320  &  Ng1543 ) ;
 assign n323 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1627) ) | ( (~ Ng853)  &  (~ Ng1621) ) | ( (~ Ng1627)  &  (~ Ng1621) ) ;
 assign n321 = ( (~ wire1594)  &  n323 ) | ( n323  &  (~ Ng1624) ) ;
 assign n325 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2081 ) | ( (~ Ng1315)  &  Ng2082 ) | ( Ng2081  &  Ng2082 ) ;
 assign n324 = ( (~ wire1603)  &  n325 ) | ( n325  &  Ng2083 ) ;
 assign n327 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2232 ) | ( (~ Ng853)  &  Ng2233 ) | ( Ng2232  &  Ng2233 ) ;
 assign n326 = ( (~ wire1594)  &  n327 ) | ( n327  &  Ng2234 ) ;
 assign n330 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2312) ) | ( (~ Ng853)  &  (~ Ng2306) ) | ( (~ Ng2312)  &  (~ Ng2306) ) ;
 assign n328 = ( (~ wire1594)  &  n330 ) | ( n330  &  (~ Ng2309) ) ;
 assign n332 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2772 ) | ( (~ Ng1315)  &  Ng2773 ) | ( Ng2772  &  Ng2773 ) ;
 assign n331 = ( (~ wire1603)  &  n332 ) | ( n332  &  Ng2774 ) ;
 assign n334 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2799 ) | ( (~ Ng1315)  &  Ng2800 ) | ( Ng2799  &  Ng2800 ) ;
 assign n333 = ( (~ wire1603)  &  n334 ) | ( n334  &  Ng2801 ) ;
 assign n337 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng192) ) | ( (~ Ng853)  &  (~ Ng186) ) | ( (~ Ng192)  &  (~ Ng186) ) ;
 assign n335 = ( (~ wire1594)  &  n337 ) | ( n337  &  (~ Ng189) ) ;
 assign n340 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng273) ) | ( (~ Ng853)  &  (~ Ng267) ) | ( (~ Ng273)  &  (~ Ng267) ) ;
 assign n338 = ( (~ wire1594)  &  n340 ) | ( n340  &  (~ Ng270) ) ;
 assign n342 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11502 ) | ( (~ Ng853)  &  Ng11500 ) | ( Ng11502  &  Ng11500 ) ;
 assign n341 = ( (~ wire1594)  &  n342 ) | ( n342  &  Ng11501 ) ;
 assign n345 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng444) ) | ( (~ Ng853)  &  (~ Ng438) ) | ( (~ Ng444)  &  (~ Ng438) ) ;
 assign n343 = ( (~ wire1594)  &  n345 ) | ( n345  &  (~ Ng441) ) ;
 assign n347 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng710 ) | ( (~ Ng1315)  &  Ng711 ) | ( Ng710  &  Ng711 ) ;
 assign n346 = ( (~ wire1603)  &  n347 ) | ( n347  &  Ng712 ) ;
 assign n349 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng820 ) | ( (~ Ng853)  &  Ng821 ) | ( Ng820  &  Ng821 ) ;
 assign n348 = ( (~ wire1594)  &  n349 ) | ( n349  &  Ng822 ) ;
 assign n352 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng951) ) | ( (~ Ng853)  &  (~ Ng945) ) | ( (~ Ng951)  &  (~ Ng945) ) ;
 assign n350 = ( (~ wire1594)  &  n352 ) | ( n352  &  (~ Ng948) ) ;
 assign n354 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11526 ) | ( (~ Ng853)  &  Ng11524 ) | ( Ng11526  &  Ng11524 ) ;
 assign n353 = ( (~ wire1594)  &  n354 ) | ( n354  &  Ng11525 ) ;
 assign n357 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1122) ) | ( (~ Ng853)  &  (~ Ng1116) ) | ( (~ Ng1122)  &  (~ Ng1116) ) ;
 assign n355 = ( (~ wire1594)  &  n357 ) | ( n357  &  (~ Ng1119) ) ;
 assign n359 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1393 ) | ( (~ Ng1315)  &  Ng1394 ) | ( Ng1393  &  Ng1394 ) ;
 assign n358 = ( (~ wire1603)  &  n359 ) | ( n359  &  Ng1395 ) ;
 assign n361 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1511 ) | ( (~ Ng853)  &  Ng1512 ) | ( Ng1511  &  Ng1512 ) ;
 assign n360 = ( (~ wire1594)  &  n361 ) | ( n361  &  Ng1513 ) ;
 assign n363 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1544 ) | ( (~ Ng853)  &  Ng1545 ) | ( Ng1544  &  Ng1545 ) ;
 assign n362 = ( (~ wire1594)  &  n363 ) | ( n363  &  Ng1546 ) ;
 assign n366 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1636) ) | ( (~ Ng853)  &  (~ Ng1630) ) | ( (~ Ng1636)  &  (~ Ng1630) ) ;
 assign n364 = ( (~ wire1594)  &  n366 ) | ( n366  &  (~ Ng1633) ) ;
 assign n368 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2084 ) | ( (~ Ng1315)  &  Ng2085 ) | ( Ng2084  &  Ng2085 ) ;
 assign n367 = ( (~ wire1603)  &  n368 ) | ( n368  &  Ng2086 ) ;
 assign n370 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2235 ) | ( (~ Ng853)  &  Ng2236 ) | ( Ng2235  &  Ng2236 ) ;
 assign n369 = ( (~ wire1594)  &  n370 ) | ( n370  &  Ng2237 ) ;
 assign n373 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2321) ) | ( (~ Ng853)  &  (~ Ng2315) ) | ( (~ Ng2321)  &  (~ Ng2315) ) ;
 assign n371 = ( (~ wire1594)  &  n373 ) | ( n373  &  (~ Ng2318) ) ;
 assign n375 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2775 ) | ( (~ Ng1315)  &  Ng2776 ) | ( Ng2775  &  Ng2776 ) ;
 assign n374 = ( (~ wire1603)  &  n375 ) | ( n375  &  Ng2777 ) ;
 assign n378 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng201) ) | ( (~ Ng853)  &  (~ Ng195) ) | ( (~ Ng201)  &  (~ Ng195) ) ;
 assign n376 = ( (~ wire1594)  &  n378 ) | ( n378  &  (~ Ng198) ) ;
 assign n380 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11505 ) | ( (~ Ng853)  &  Ng11503 ) | ( Ng11505  &  Ng11503 ) ;
 assign n379 = ( (~ wire1594)  &  n380 ) | ( n380  &  Ng11504 ) ;
 assign n382 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng713 ) | ( (~ Ng1315)  &  Ng714 ) | ( Ng713  &  Ng714 ) ;
 assign n381 = ( (~ wire1603)  &  n382 ) | ( n382  &  Ng715 ) ;
 assign n384 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng731 ) | ( (~ Ng1315)  &  Ng732 ) | ( Ng731  &  Ng732 ) ;
 assign n383 = ( (~ wire1603)  &  n384 ) | ( n384  &  Ng733 ) ;
 assign n387 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng879) ) | ( (~ Ng853)  &  (~ Ng873) ) | ( (~ Ng879)  &  (~ Ng873) ) ;
 assign n385 = ( (~ wire1594)  &  n387 ) | ( n387  &  (~ Ng876) ) ;
 assign n390 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng960) ) | ( (~ Ng853)  &  (~ Ng954) ) | ( (~ Ng960)  &  (~ Ng954) ) ;
 assign n388 = ( (~ wire1594)  &  n390 ) | ( n390  &  (~ Ng957) ) ;
 assign n392 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11529 ) | ( (~ Ng853)  &  Ng11527 ) | ( Ng11529  &  Ng11527 ) ;
 assign n391 = ( (~ wire1594)  &  n392 ) | ( n392  &  Ng11528 ) ;
 assign n395 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1131) ) | ( (~ Ng853)  &  (~ Ng1125) ) | ( (~ Ng1131)  &  (~ Ng1125) ) ;
 assign n393 = ( (~ wire1594)  &  n395 ) | ( n395  &  (~ Ng1128) ) ;
 assign n397 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1396 ) | ( (~ Ng1315)  &  Ng1397 ) | ( Ng1396  &  Ng1397 ) ;
 assign n396 = ( (~ wire1603)  &  n397 ) | ( n397  &  Ng1398 ) ;
 assign n399 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1514 ) | ( (~ Ng853)  &  Ng1515 ) | ( Ng1514  &  Ng1515 ) ;
 assign n398 = ( (~ wire1594)  &  n399 ) | ( n399  &  Ng1516 ) ;
 assign n402 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1645) ) | ( (~ Ng853)  &  (~ Ng1639) ) | ( (~ Ng1645)  &  (~ Ng1639) ) ;
 assign n400 = ( (~ wire1594)  &  n402 ) | ( n402  &  (~ Ng1642) ) ;
 assign n404 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11553 ) | ( (~ Ng853)  &  Ng11551 ) | ( Ng11553  &  Ng11551 ) ;
 assign n403 = ( (~ wire1594)  &  n404 ) | ( n404  &  Ng11552 ) ;
 assign n407 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1816) ) | ( (~ Ng853)  &  (~ Ng1810) ) | ( (~ Ng1816)  &  (~ Ng1810) ) ;
 assign n405 = ( (~ wire1594)  &  n407 ) | ( n407  &  (~ Ng1813) ) ;
 assign n409 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2087 ) | ( (~ Ng1315)  &  Ng2088 ) | ( Ng2087  &  Ng2088 ) ;
 assign n408 = ( (~ wire1603)  &  n409 ) | ( n409  &  Ng2089 ) ;
 assign n411 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2205 ) | ( (~ Ng853)  &  Ng2206 ) | ( Ng2205  &  Ng2206 ) ;
 assign n410 = ( (~ wire1594)  &  n411 ) | ( n411  &  Ng2207 ) ;
 assign n413 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2238 ) | ( (~ Ng853)  &  Ng2239 ) | ( Ng2238  &  Ng2239 ) ;
 assign n412 = ( (~ wire1594)  &  n413 ) | ( n413  &  Ng2240 ) ;
 assign n416 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2330) ) | ( (~ Ng853)  &  (~ Ng2324) ) | ( (~ Ng2330)  &  (~ Ng2324) ) ;
 assign n414 = ( (~ wire1594)  &  n416 ) | ( n416  &  (~ Ng2327) ) ;
 assign n418 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2778 ) | ( (~ Ng1315)  &  Ng2779 ) | ( Ng2778  &  Ng2779 ) ;
 assign n417 = ( (~ wire1603)  &  n418 ) | ( n418  &  Ng2780 ) ;
 assign n421 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng210) ) | ( (~ Ng853)  &  (~ Ng204) ) | ( (~ Ng210)  &  (~ Ng204) ) ;
 assign n419 = ( (~ wire1594)  &  n421 ) | ( n421  &  (~ Ng207) ) ;
 assign n423 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11508 ) | ( (~ Ng853)  &  Ng11506 ) | ( Ng11508  &  Ng11506 ) ;
 assign n422 = ( (~ wire1594)  &  n423 ) | ( n423  &  Ng11507 ) ;
 assign n425 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng716 ) | ( (~ Ng1315)  &  Ng717 ) | ( Ng716  &  Ng717 ) ;
 assign n424 = ( (~ wire1603)  &  n425 ) | ( n425  &  Ng718 ) ;
 assign n428 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng888) ) | ( (~ Ng853)  &  (~ Ng882) ) | ( (~ Ng888)  &  (~ Ng882) ) ;
 assign n426 = ( (~ wire1594)  &  n428 ) | ( n428  &  (~ Ng885) ) ;
 assign n430 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11532 ) | ( (~ Ng853)  &  Ng11530 ) | ( Ng11532  &  Ng11530 ) ;
 assign n429 = ( (~ wire1594)  &  n430 ) | ( n430  &  Ng11531 ) ;
 assign n432 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1399 ) | ( (~ Ng1315)  &  Ng1400 ) | ( Ng1399  &  Ng1400 ) ;
 assign n431 = ( (~ wire1603)  &  n432 ) | ( n432  &  Ng1401 ) ;
 assign n434 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1417 ) | ( (~ Ng1315)  &  Ng1418 ) | ( Ng1417  &  Ng1418 ) ;
 assign n433 = ( (~ wire1603)  &  n434 ) | ( n434  &  Ng1419 ) ;
 assign n437 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1573) ) | ( (~ Ng853)  &  (~ Ng1567) ) | ( (~ Ng1573)  &  (~ Ng1567) ) ;
 assign n435 = ( (~ wire1594)  &  n437 ) | ( n437  &  (~ Ng1570) ) ;
 assign n440 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1654) ) | ( (~ Ng853)  &  (~ Ng1648) ) | ( (~ Ng1654)  &  (~ Ng1648) ) ;
 assign n438 = ( (~ wire1594)  &  n440 ) | ( n440  &  (~ Ng1651) ) ;
 assign n442 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11556 ) | ( (~ Ng853)  &  Ng11554 ) | ( Ng11556  &  Ng11554 ) ;
 assign n441 = ( (~ wire1594)  &  n442 ) | ( n442  &  Ng11555 ) ;
 assign n445 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1825) ) | ( (~ Ng853)  &  (~ Ng1819) ) | ( (~ Ng1825)  &  (~ Ng1819) ) ;
 assign n443 = ( (~ wire1594)  &  n445 ) | ( n445  &  (~ Ng1822) ) ;
 assign n447 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2090 ) | ( (~ Ng1315)  &  Ng2091 ) | ( Ng2090  &  Ng2091 ) ;
 assign n446 = ( (~ wire1603)  &  n447 ) | ( n447  &  Ng2092 ) ;
 assign n449 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2208 ) | ( (~ Ng853)  &  Ng2209 ) | ( Ng2208  &  Ng2209 ) ;
 assign n448 = ( (~ wire1594)  &  n449 ) | ( n449  &  Ng2210 ) ;
 assign n452 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2339) ) | ( (~ Ng853)  &  (~ Ng2333) ) | ( (~ Ng2339)  &  (~ Ng2333) ) ;
 assign n450 = ( (~ wire1594)  &  n452 ) | ( n452  &  (~ Ng2336) ) ;
 assign n454 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11580 ) | ( (~ Ng853)  &  Ng11578 ) | ( Ng11580  &  Ng11578 ) ;
 assign n453 = ( (~ wire1594)  &  n454 ) | ( n454  &  Ng11579 ) ;
 assign n457 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2510) ) | ( (~ Ng853)  &  (~ Ng2504) ) | ( (~ Ng2510)  &  (~ Ng2504) ) ;
 assign n455 = ( (~ wire1594)  &  n457 ) | ( n457  &  (~ Ng2507) ) ;
 assign n459 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2781 ) | ( (~ Ng1315)  &  Ng2782 ) | ( Ng2781  &  Ng2782 ) ;
 assign n458 = ( (~ wire1603)  &  n459 ) | ( n459  &  Ng2783 ) ;
 assign n461 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng168 ) | ( (~ Ng853)  &  Ng170 ) | ( Ng168  &  Ng170 ) ;
 assign n460 = ( (~ wire1612)  &  n461 ) | ( n461  &  Ng169 ) ;
 assign n463 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng719 ) | ( (~ Ng1315)  &  Ng720 ) | ( Ng719  &  Ng720 ) ;
 assign n462 = ( (~ wire1603)  &  n463 ) | ( n463  &  Ng721 ) ;
 assign n466 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng897) ) | ( (~ Ng853)  &  (~ Ng891) ) | ( (~ Ng897)  &  (~ Ng891) ) ;
 assign n464 = ( (~ wire1594)  &  n466 ) | ( n466  &  (~ Ng894) ) ;
 assign n468 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11535 ) | ( (~ Ng853)  &  Ng11533 ) | ( Ng11535  &  Ng11533 ) ;
 assign n467 = ( (~ wire1594)  &  n468 ) | ( n468  &  Ng11534 ) ;
 assign n470 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1402 ) | ( (~ Ng1315)  &  Ng1403 ) | ( Ng1402  &  Ng1403 ) ;
 assign n469 = ( (~ wire1603)  &  n470 ) | ( n470  &  Ng1404 ) ;
 assign n473 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1582) ) | ( (~ Ng853)  &  (~ Ng1576) ) | ( (~ Ng1582)  &  (~ Ng1576) ) ;
 assign n471 = ( (~ wire1594)  &  n473 ) | ( n473  &  (~ Ng1579) ) ;
 assign n475 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11559 ) | ( (~ Ng853)  &  Ng11557 ) | ( Ng11559  &  Ng11557 ) ;
 assign n474 = ( (~ wire1594)  &  n475 ) | ( n475  &  Ng11558 ) ;
 assign n477 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2093 ) | ( (~ Ng1315)  &  Ng2094 ) | ( Ng2093  &  Ng2094 ) ;
 assign n476 = ( (~ wire1603)  &  n477 ) | ( n477  &  Ng2095 ) ;
 assign n479 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2111 ) | ( (~ Ng1315)  &  Ng2112 ) | ( Ng2111  &  Ng2112 ) ;
 assign n478 = ( (~ wire1603)  &  n479 ) | ( n479  &  Ng2113 ) ;
 assign n482 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2267) ) | ( (~ Ng853)  &  (~ Ng2261) ) | ( (~ Ng2267)  &  (~ Ng2261) ) ;
 assign n480 = ( (~ wire1594)  &  n482 ) | ( n482  &  (~ Ng2264) ) ;
 assign n485 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2348) ) | ( (~ Ng853)  &  (~ Ng2342) ) | ( (~ Ng2348)  &  (~ Ng2342) ) ;
 assign n483 = ( (~ wire1594)  &  n485 ) | ( n485  &  (~ Ng2345) ) ;
 assign n487 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11583 ) | ( (~ Ng853)  &  Ng11581 ) | ( Ng11583  &  Ng11581 ) ;
 assign n486 = ( (~ wire1594)  &  n487 ) | ( n487  &  Ng11582 ) ;
 assign n490 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2519) ) | ( (~ Ng853)  &  (~ Ng2513) ) | ( (~ Ng2519)  &  (~ Ng2513) ) ;
 assign n488 = ( (~ wire1594)  &  n490 ) | ( n490  &  (~ Ng2516) ) ;
 assign n492 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2784 ) | ( (~ Ng1315)  &  Ng2785 ) | ( Ng2784  &  Ng2785 ) ;
 assign n491 = ( (~ wire1603)  &  n492 ) | ( n492  &  Ng2786 ) ;
 assign n494 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng722 ) | ( (~ Ng1315)  &  Ng723 ) | ( Ng722  &  Ng723 ) ;
 assign n493 = ( (~ wire1603)  &  n494 ) | ( n494  &  Ng724 ) ;
 assign n496 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng856 ) | ( (~ Ng853)  &  Ng858 ) | ( Ng856  &  Ng858 ) ;
 assign n495 = ( (~ wire1612)  &  n496 ) | ( n496  &  Ng857 ) ;
 assign n498 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1405 ) | ( (~ Ng1315)  &  Ng1406 ) | ( Ng1405  &  Ng1406 ) ;
 assign n497 = ( (~ wire1603)  &  n498 ) | ( n498  &  Ng1407 ) ;
 assign n501 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1591) ) | ( (~ Ng853)  &  (~ Ng1585) ) | ( (~ Ng1591)  &  (~ Ng1585) ) ;
 assign n499 = ( (~ wire1594)  &  n501 ) | ( n501  &  (~ Ng1588) ) ;
 assign n503 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11562 ) | ( (~ Ng853)  &  Ng11560 ) | ( Ng11562  &  Ng11560 ) ;
 assign n502 = ( (~ wire1594)  &  n503 ) | ( n503  &  Ng11561 ) ;
 assign n505 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2096 ) | ( (~ Ng1315)  &  Ng2097 ) | ( Ng2096  &  Ng2097 ) ;
 assign n504 = ( (~ wire1603)  &  n505 ) | ( n505  &  Ng2098 ) ;
 assign n508 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2276) ) | ( (~ Ng853)  &  (~ Ng2270) ) | ( (~ Ng2276)  &  (~ Ng2270) ) ;
 assign n506 = ( (~ wire1594)  &  n508 ) | ( n508  &  (~ Ng2273) ) ;
 assign n510 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11586 ) | ( (~ Ng853)  &  Ng11584 ) | ( Ng11586  &  Ng11584 ) ;
 assign n509 = ( (~ wire1594)  &  n510 ) | ( n510  &  Ng11585 ) ;
 assign n512 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2787 ) | ( (~ Ng1315)  &  Ng2788 ) | ( Ng2787  &  Ng2788 ) ;
 assign n511 = ( (~ wire1603)  &  n512 ) | ( n512  &  Ng2789 ) ;
 assign n514 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2805 ) | ( (~ Ng1315)  &  Ng2806 ) | ( Ng2805  &  Ng2806 ) ;
 assign n513 = ( (~ wire1603)  &  n514 ) | ( n514  &  Ng2807 ) ;
 assign n516 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1408 ) | ( (~ Ng1315)  &  Ng1409 ) | ( Ng1408  &  Ng1409 ) ;
 assign n515 = ( (~ wire1603)  &  n516 ) | ( n516  &  Ng1410 ) ;
 assign n518 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1550 ) | ( (~ Ng853)  &  Ng1551 ) | ( Ng1550  &  Ng1551 ) ;
 assign n517 = ( (~ wire1594)  &  n518 ) | ( n518  &  Ng1552 ) ;
 assign n520 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2099 ) | ( (~ Ng1315)  &  Ng2100 ) | ( Ng2099  &  Ng2100 ) ;
 assign n519 = ( (~ wire1603)  &  n520 ) | ( n520  &  Ng2101 ) ;
 assign n523 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2285) ) | ( (~ Ng853)  &  (~ Ng2279) ) | ( (~ Ng2285)  &  (~ Ng2279) ) ;
 assign n521 = ( (~ wire1594)  &  n523 ) | ( n523  &  (~ Ng2282) ) ;
 assign n525 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng11589 ) | ( (~ Ng853)  &  Ng11587 ) | ( Ng11589  &  Ng11587 ) ;
 assign n524 = ( (~ wire1594)  &  n525 ) | ( n525  &  Ng11588 ) ;
 assign n527 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2790 ) | ( (~ Ng1315)  &  Ng2791 ) | ( Ng2790  &  Ng2791 ) ;
 assign n526 = ( (~ wire1603)  &  n527 ) | ( n527  &  Ng2792 ) ;
 assign n529 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2102 ) | ( (~ Ng1315)  &  Ng2103 ) | ( Ng2102  &  Ng2103 ) ;
 assign n528 = ( (~ wire1603)  &  n529 ) | ( n529  &  Ng2104 ) ;
 assign n531 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2244 ) | ( (~ Ng853)  &  Ng2245 ) | ( Ng2244  &  Ng2245 ) ;
 assign n530 = ( (~ wire1594)  &  n531 ) | ( n531  &  Ng2246 ) ;
 assign n533 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2793 ) | ( (~ Ng1315)  &  Ng2794 ) | ( Ng2793  &  Ng2794 ) ;
 assign n532 = ( (~ wire1603)  &  n533 ) | ( n533  &  Ng2795 ) ;
 assign n535 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng314 ) | ( (~ Ng853)  &  Ng312 ) | ( Ng314  &  Ng312 ) ;
 assign n534 = ( (~ wire1594)  &  n535 ) | ( n535  &  Ng313 ) ;
 assign n537 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2796 ) | ( (~ Ng1315)  &  Ng2797 ) | ( Ng2796  &  Ng2797 ) ;
 assign n536 = ( (~ wire1603)  &  n537 ) | ( n537  &  Ng2798 ) ;
 assign n539 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng317 ) | ( (~ Ng853)  &  Ng315 ) | ( Ng317  &  Ng315 ) ;
 assign n538 = ( (~ wire1594)  &  n539 ) | ( n539  &  Ng316 ) ;
 assign n541 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1001 ) | ( (~ Ng853)  &  Ng999 ) | ( Ng1001  &  Ng999 ) ;
 assign n540 = ( (~ wire1594)  &  n541 ) | ( n541  &  Ng1000 ) ;
 assign n543 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng320 ) | ( (~ Ng853)  &  Ng318 ) | ( Ng320  &  Ng318 ) ;
 assign n542 = ( (~ wire1594)  &  n543 ) | ( n543  &  Ng319 ) ;
 assign n545 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1004 ) | ( (~ Ng853)  &  Ng1002 ) | ( Ng1004  &  Ng1002 ) ;
 assign n544 = ( (~ wire1594)  &  n545 ) | ( n545  &  Ng1003 ) ;
 assign n547 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1695 ) | ( (~ Ng853)  &  Ng1693 ) | ( Ng1695  &  Ng1693 ) ;
 assign n546 = ( (~ wire1594)  &  n547 ) | ( n547  &  Ng1694 ) ;
 assign n550 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng620) ) | ( (~ Ng1315)  &  (~ Ng614) ) | ( (~ Ng620)  &  (~ Ng614) ) ;
 assign n548 = ( (~ wire1603)  &  n550 ) | ( n550  &  (~ Ng617) ) ;
 assign n552 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1007 ) | ( (~ Ng853)  &  Ng1005 ) | ( Ng1007  &  Ng1005 ) ;
 assign n551 = ( (~ wire1594)  &  n552 ) | ( n552  &  Ng1006 ) ;
 assign n554 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1698 ) | ( (~ Ng853)  &  Ng1696 ) | ( Ng1698  &  Ng1696 ) ;
 assign n553 = ( (~ wire1594)  &  n554 ) | ( n554  &  Ng1697 ) ;
 assign n556 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2389 ) | ( (~ Ng853)  &  Ng2387 ) | ( Ng2389  &  Ng2387 ) ;
 assign n555 = ( (~ wire1594)  &  n556 ) | ( n556  &  Ng2388 ) ;
 assign n559 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1306) ) | ( (~ Ng1315)  &  (~ Ng1300) ) | ( (~ Ng1306)  &  (~ Ng1300) ) ;
 assign n557 = ( (~ wire1603)  &  n559 ) | ( n559  &  (~ Ng1303) ) ;
 assign n561 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1701 ) | ( (~ Ng853)  &  Ng1699 ) | ( Ng1701  &  Ng1699 ) ;
 assign n560 = ( (~ wire1594)  &  n561 ) | ( n561  &  Ng1700 ) ;
 assign n563 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2392 ) | ( (~ Ng853)  &  Ng2390 ) | ( Ng2392  &  Ng2390 ) ;
 assign n562 = ( (~ wire1594)  &  n563 ) | ( n563  &  Ng2391 ) ;
 assign n566 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2000) ) | ( (~ Ng1315)  &  (~ Ng1994) ) | ( (~ Ng2000)  &  (~ Ng1994) ) ;
 assign n564 = ( (~ wire1603)  &  n566 ) | ( n566  &  (~ Ng1997) ) ;
 assign n568 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2395 ) | ( (~ Ng853)  &  Ng2393 ) | ( Ng2395  &  Ng2393 ) ;
 assign n567 = ( (~ wire1594)  &  n568 ) | ( n568  &  Ng2394 ) ;
 assign n571 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2694) ) | ( (~ Ng1315)  &  (~ Ng2688) ) | ( (~ Ng2694)  &  (~ Ng2688) ) ;
 assign n569 = ( (~ wire1603)  &  n571 ) | ( n571  &  (~ Ng2691) ) ;
 assign n573 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng575 ) | ( (~ Ng1315)  &  Ng576 ) | ( Ng575  &  Ng576 ) ;
 assign n572 = ( (~ wire1603)  &  n573 ) | ( n573  &  Ng577 ) ;
 assign n575 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng578 ) | ( (~ Ng1315)  &  Ng579 ) | ( Ng578  &  Ng579 ) ;
 assign n574 = ( (~ wire1603)  &  n575 ) | ( n575  &  Ng580 ) ;
 assign n577 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1261 ) | ( (~ Ng1315)  &  Ng1262 ) | ( Ng1261  &  Ng1262 ) ;
 assign n576 = ( (~ wire1603)  &  n577 ) | ( n577  &  Ng1263 ) ;
 assign n580 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng414) ) | ( (~ Ng853)  &  (~ Ng408) ) | ( (~ Ng414)  &  (~ Ng408) ) ;
 assign n578 = ( (~ wire1594)  &  n580 ) | ( n580  &  (~ Ng411) ) ;
 assign n582 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng581 ) | ( (~ Ng1315)  &  Ng582 ) | ( Ng581  &  Ng582 ) ;
 assign n581 = ( (~ wire1603)  &  n582 ) | ( n582  &  Ng583 ) ;
 assign n584 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1264 ) | ( (~ Ng1315)  &  Ng1265 ) | ( Ng1264  &  Ng1265 ) ;
 assign n583 = ( (~ wire1603)  &  n584 ) | ( n584  &  Ng1266 ) ;
 assign n586 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1955 ) | ( (~ Ng1315)  &  Ng1956 ) | ( Ng1955  &  Ng1956 ) ;
 assign n585 = ( (~ wire1603)  &  n586 ) | ( n586  &  Ng1957 ) ;
 assign n589 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng423) ) | ( (~ Ng853)  &  (~ Ng417) ) | ( (~ Ng423)  &  (~ Ng417) ) ;
 assign n587 = ( (~ wire1594)  &  n589 ) | ( n589  &  (~ Ng420) ) ;
 assign n591 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng584 ) | ( (~ Ng1315)  &  Ng585 ) | ( Ng584  &  Ng585 ) ;
 assign n590 = ( (~ wire1603)  &  n591 ) | ( n591  &  Ng586 ) ;
 assign n594 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1101) ) | ( (~ Ng853)  &  (~ Ng1095) ) | ( (~ Ng1101)  &  (~ Ng1095) ) ;
 assign n592 = ( (~ wire1594)  &  n594 ) | ( n594  &  (~ Ng1098) ) ;
 assign n596 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1267 ) | ( (~ Ng1315)  &  Ng1268 ) | ( Ng1267  &  Ng1268 ) ;
 assign n595 = ( (~ wire1603)  &  n596 ) | ( n596  &  Ng1269 ) ;
 assign n598 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1958 ) | ( (~ Ng1315)  &  Ng1959 ) | ( Ng1958  &  Ng1959 ) ;
 assign n597 = ( (~ wire1603)  &  n598 ) | ( n598  &  Ng1960 ) ;
 assign n600 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2649 ) | ( (~ Ng1315)  &  Ng2650 ) | ( Ng2649  &  Ng2650 ) ;
 assign n599 = ( (~ wire1603)  &  n600 ) | ( n600  &  Ng2651 ) ;
 assign n603 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1110) ) | ( (~ Ng853)  &  (~ Ng1104) ) | ( (~ Ng1110)  &  (~ Ng1104) ) ;
 assign n601 = ( (~ wire1594)  &  n603 ) | ( n603  &  (~ Ng1107) ) ;
 assign n605 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1270 ) | ( (~ Ng1315)  &  Ng1271 ) | ( Ng1270  &  Ng1271 ) ;
 assign n604 = ( (~ wire1603)  &  n605 ) | ( n605  &  Ng1272 ) ;
 assign n608 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1795) ) | ( (~ Ng853)  &  (~ Ng1789) ) | ( (~ Ng1795)  &  (~ Ng1789) ) ;
 assign n606 = ( (~ wire1594)  &  n608 ) | ( n608  &  (~ Ng1792) ) ;
 assign n610 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1961 ) | ( (~ Ng1315)  &  Ng1962 ) | ( Ng1961  &  Ng1962 ) ;
 assign n609 = ( (~ wire1603)  &  n610 ) | ( n610  &  Ng1963 ) ;
 assign n612 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2652 ) | ( (~ Ng1315)  &  Ng2653 ) | ( Ng2652  &  Ng2653 ) ;
 assign n611 = ( (~ wire1603)  &  n612 ) | ( n612  &  Ng2654 ) ;
 assign n614 = ( (~ wire1594)  &  (~ Ng853) ) | ( (~ wire1594)  &  Ng171 ) | ( (~ Ng853)  &  Ng173 ) | ( Ng171  &  Ng173 ) ;
 assign n613 = ( (~ wire1612)  &  n614 ) | ( n614  &  Ng172 ) ;
 assign n617 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng1804) ) | ( (~ Ng853)  &  (~ Ng1798) ) | ( (~ Ng1804)  &  (~ Ng1798) ) ;
 assign n615 = ( (~ wire1594)  &  n617 ) | ( n617  &  (~ Ng1801) ) ;
 assign n619 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng1964 ) | ( (~ Ng1315)  &  Ng1965 ) | ( Ng1964  &  Ng1965 ) ;
 assign n618 = ( (~ wire1603)  &  n619 ) | ( n619  &  Ng1966 ) ;
 assign n622 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2489) ) | ( (~ Ng853)  &  (~ Ng2483) ) | ( (~ Ng2489)  &  (~ Ng2483) ) ;
 assign n620 = ( (~ wire1594)  &  n622 ) | ( n622  &  (~ Ng2486) ) ;
 assign n624 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2655 ) | ( (~ Ng1315)  &  Ng2656 ) | ( Ng2655  &  Ng2656 ) ;
 assign n623 = ( (~ wire1603)  &  n624 ) | ( n624  &  Ng2657 ) ;
 assign n626 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng174 ) | ( (~ Ng853)  &  Ng175 ) | ( Ng174  &  Ng175 ) ;
 assign n625 = ( (~ wire1594)  &  n626 ) | ( n626  &  Ng176 ) ;
 assign n628 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng859 ) | ( (~ Ng853)  &  Ng860 ) | ( Ng859  &  Ng860 ) ;
 assign n627 = ( (~ wire1594)  &  n628 ) | ( n628  &  Ng861 ) ;
 assign n631 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  (~ Ng2498) ) | ( (~ Ng853)  &  (~ Ng2492) ) | ( (~ Ng2498)  &  (~ Ng2492) ) ;
 assign n629 = ( (~ wire1594)  &  n631 ) | ( n631  &  (~ Ng2495) ) ;
 assign n633 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  Ng2658 ) | ( (~ Ng1315)  &  Ng2659 ) | ( Ng2658  &  Ng2659 ) ;
 assign n632 = ( (~ wire1603)  &  n633 ) | ( n633  &  Ng2660 ) ;
 assign n635 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng862 ) | ( (~ Ng853)  &  Ng863 ) | ( Ng862  &  Ng863 ) ;
 assign n634 = ( (~ wire1594)  &  n635 ) | ( n635  &  Ng864 ) ;
 assign n637 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1553 ) | ( (~ Ng853)  &  Ng1554 ) | ( Ng1553  &  Ng1554 ) ;
 assign n636 = ( (~ wire1594)  &  n637 ) | ( n637  &  Ng1555 ) ;
 assign n639 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1556 ) | ( (~ Ng853)  &  Ng1557 ) | ( Ng1556  &  Ng1557 ) ;
 assign n638 = ( (~ wire1594)  &  n639 ) | ( n639  &  Ng1558 ) ;
 assign n641 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2247 ) | ( (~ Ng853)  &  Ng2248 ) | ( Ng2247  &  Ng2248 ) ;
 assign n640 = ( (~ wire1594)  &  n641 ) | ( n641  &  Ng2249 ) ;
 assign n643 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2250 ) | ( (~ Ng853)  &  Ng2251 ) | ( Ng2250  &  Ng2251 ) ;
 assign n642 = ( (~ wire1594)  &  n643 ) | ( n643  &  Ng2252 ) ;
 assign n644 = ( (~ Pg8021)  &  Ng2879 ) | ( Ng2879  &  Ng2929 ) ;
 assign Ng16494 = ( (~ n644) ) ;
 assign n646 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ Ng853)  &  Ng427 ) | ( (~ wire1612)  &  Ng426 ) | ( Ng427  &  Ng426 ) ;
 assign n645 = ( (~ wire1594)  &  n646 ) | ( n646  &  Ng428 ) ;
 assign n648 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ Ng853)  &  Ng1114 ) | ( (~ wire1612)  &  Ng1113 ) | ( Ng1114  &  Ng1113 ) ;
 assign n647 = ( (~ wire1594)  &  n648 ) | ( n648  &  Ng1115 ) ;
 assign n651 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng611) ) | ( (~ Ng1315)  &  (~ Ng605) ) | ( (~ Ng611)  &  (~ Ng605) ) ;
 assign n649 = ( (~ wire1603)  &  n651 ) | ( n651  &  (~ Ng608) ) ;
 assign n653 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ Ng853)  &  Ng1808 ) | ( (~ wire1612)  &  Ng1807 ) | ( Ng1808  &  Ng1807 ) ;
 assign n652 = ( (~ wire1594)  &  n653 ) | ( n653  &  Ng1809 ) ;
 assign n656 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1297) ) | ( (~ Ng1315)  &  (~ Ng1291) ) | ( (~ Ng1297)  &  (~ Ng1291) ) ;
 assign n654 = ( (~ wire1603)  &  n656 ) | ( n656  &  (~ Ng1294) ) ;
 assign n658 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ Ng853)  &  Ng2502 ) | ( (~ wire1612)  &  Ng2501 ) | ( Ng2502  &  Ng2501 ) ;
 assign n657 = ( (~ wire1594)  &  n658 ) | ( n658  &  Ng2503 ) ;
 assign n661 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1991) ) | ( (~ Ng1315)  &  (~ Ng1985) ) | ( (~ Ng1991)  &  (~ Ng1985) ) ;
 assign n659 = ( (~ wire1603)  &  n661 ) | ( n661  &  (~ Ng1988) ) ;
 assign n664 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2685) ) | ( (~ Ng1315)  &  (~ Ng2679) ) | ( (~ Ng2685)  &  (~ Ng2679) ) ;
 assign n662 = ( (~ wire1603)  &  n664 ) | ( n664  &  (~ Ng2682) ) ;
 assign n665 = ( Ng525  &  (~ Ng557) ) | ( Ng510  &  (~ Ng557) ) ;
 assign n667 = ( Ng525  &  (~ Ng510) ) | ( (~ Ng510)  &  Ng557 ) ;
 assign n669 = ( Ng1211  &  (~ Ng1243) ) | ( Ng1196  &  (~ Ng1243) ) ;
 assign n671 = ( Ng1211  &  (~ Ng1196) ) | ( (~ Ng1196)  &  Ng1243 ) ;
 assign n673 = ( Ng1905  &  (~ Ng1937) ) | ( Ng1890  &  (~ Ng1937) ) ;
 assign n675 = ( Ng1905  &  (~ Ng1890) ) | ( (~ Ng1890)  &  Ng1937 ) ;
 assign n677 = ( Ng2599  &  (~ Ng2631) ) | ( Ng2584  &  (~ Ng2631) ) ;
 assign n679 = ( Ng2599  &  (~ Ng2584) ) | ( (~ Ng2584)  &  Ng2631 ) ;
 assign n683 = ( Ng16467 ) | ( (~ Ng185) ) | ( (~ Ng524) ) ;
 assign n684 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng593) ) | ( (~ Ng1315)  &  (~ Ng587) ) | ( (~ Ng593)  &  (~ Ng587) ) ;
 assign n681 = ( (~ wire1603)  &  n683  &  n684 ) | ( n683  &  n684  &  (~ Ng590) ) ;
 assign n687 = ( Ng16469 ) | ( (~ Ng185) ) | ( (~ Ng1210) ) ;
 assign n688 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1279) ) | ( (~ Ng1315)  &  (~ Ng1273) ) | ( (~ Ng1279)  &  (~ Ng1273) ) ;
 assign n685 = ( (~ wire1603)  &  n687  &  n688 ) | ( n687  &  n688  &  (~ Ng1276) ) ;
 assign n691 = ( Ng16471 ) | ( (~ Ng185) ) | ( (~ Ng1904) ) ;
 assign n692 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng1973) ) | ( (~ Ng1315)  &  (~ Ng1967) ) | ( (~ Ng1973)  &  (~ Ng1967) ) ;
 assign n689 = ( (~ wire1603)  &  n691  &  n692 ) | ( n691  &  n692  &  (~ Ng1970) ) ;
 assign n695 = ( Ng16473 ) | ( (~ Ng185) ) | ( (~ Ng2598) ) ;
 assign n696 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ wire1605)  &  (~ Ng2667) ) | ( (~ Ng1315)  &  (~ Ng2661) ) | ( (~ Ng2667)  &  (~ Ng2661) ) ;
 assign n693 = ( (~ wire1603)  &  n695  &  n696 ) | ( n695  &  n696  &  (~ Ng2664) ) ;
 assign Ng20571 = ( (~ Pg51)  &  Ng13457 ) ;
 assign Ng20588 = ( (~ Pg51)  &  Ng2817 ) ;
 assign n698 = ( (~ Ng659)  &  n1960 ) | ( n1960  &  n1958 ) ;
 assign Ng21943 = ( (~ n698) ) ;
 assign n699 = ( (~ Ng1345)  &  n1960 ) | ( n1960  &  n1958 ) ;
 assign Ng21944 = ( (~ n699) ) ;
 assign n700 = ( (~ Ng2039)  &  n1960 ) | ( n1960  &  n1958 ) ;
 assign Ng21945 = ( (~ n700) ) ;
 assign n701 = ( (~ Ng2733)  &  n1960 ) | ( n1960  &  n1958 ) ;
 assign Ng21946 = ( (~ n701) ) ;
 assign Ng21951 = ( Pg51 ) | ( Ng2933 ) ;
 assign Ng21965 = ( Ng3079 ) | ( Pg3234 ) ;
 assign n702 = ( n1951  &  n1949 ) | ( n1951  &  (~ Ng554) ) ;
 assign Ng23160 = ( (~ n702) ) ;
 assign n703 = ( n1951  &  n1949 ) | ( n1951  &  (~ Ng1240) ) ;
 assign Ng23198 = ( (~ n703) ) ;
 assign n704 = ( n1951  &  n1949 ) | ( n1951  &  (~ Ng1934) ) ;
 assign Ng23236 = ( (~ n704) ) ;
 assign n705 = ( n1951  &  n1949 ) | ( n1951  &  (~ Ng2628) ) ;
 assign Ng23274 = ( (~ n705) ) ;
 assign n706 = ( n1956  &  Ng640 ) | ( (~ n1956)  &  (~ Ng640) ) ;
 assign n707 = ( (~ wire1603) ) | ( (~ Ng630) ) ;
 assign Ng23161 = ( n706  &  n707 ) ;
 assign n708 = ( n1954  &  Ng1326 ) | ( (~ n1954)  &  (~ Ng1326) ) ;
 assign n709 = ( (~ wire1603) ) | ( (~ Ng1316) ) ;
 assign Ng23199 = ( n708  &  n709 ) ;
 assign n710 = ( n1952  &  Ng2020 ) | ( (~ n1952)  &  (~ Ng2020) ) ;
 assign n711 = ( (~ wire1603) ) | ( (~ Ng2010) ) ;
 assign Ng23237 = ( n710  &  n711 ) ;
 assign n712 = ( n1948  &  Ng2714 ) | ( (~ n1948)  &  (~ Ng2714) ) ;
 assign n713 = ( (~ wire1603) ) | ( (~ Ng2704) ) ;
 assign Ng23275 = ( n712  &  n713 ) ;
 assign n714 = ( n1938 ) | ( Pg8021 ) ;
 assign n715 = ( (~ Ng2883)  &  Ng13457 ) | ( Ng2883  &  (~ Ng13457) ) ;
 assign Ng23315 = ( n714 ) | ( n715 ) ;
 assign Ng23317 = ( (~ Pg3234)  &  Ng13475 ) ;
 assign Ng23318 = ( (~ Pg3234)  &  Ng3054 ) ;
 assign n717 = ( (~ n1946)  &  Ng633 ) | ( n1946  &  (~ Ng633) ) ;
 assign Ng24296 = ( n717  &  n707 ) ;
 assign n718 = ( (~ n1944)  &  Ng1319 ) | ( n1944  &  (~ Ng1319) ) ;
 assign Ng24337 = ( n718  &  n709 ) ;
 assign n722 = ( (~ n534) ) | ( n538 ) | ( n542 ) ;
 assign n721 = ( Ng2892 ) | ( Ng2903 ) | ( Ng2908 ) | ( Ng2896 ) | ( Ng2900 ) ;
 assign n719 = ( n722  &  n721 ) | ( n722  &  (~ n1901) ) ;
 assign n723 = ( (~ n1942)  &  Ng2013 ) | ( n1942  &  (~ Ng2013) ) ;
 assign Ng24378 = ( n723  &  n711 ) ;
 assign n726 = ( (~ n540) ) | ( n544 ) | ( n551 ) ;
 assign n724 = ( n721  &  n726 ) | ( n726  &  (~ n1897) ) ;
 assign n727 = ( (~ n1940)  &  Ng2707 ) | ( n1940  &  (~ Ng2707) ) ;
 assign Ng24419 = ( n727  &  n713 ) ;
 assign n730 = ( (~ n546) ) | ( n553 ) | ( n560 ) ;
 assign n728 = ( n721  &  n730 ) | ( n730  &  (~ n1893) ) ;
 assign n733 = ( (~ n555) ) | ( n562 ) | ( n567 ) ;
 assign n731 = ( n721  &  n733 ) | ( n733  &  (~ n1889) ) ;
 assign n734 = ( n714  &  Pg8021 ) | ( n714  &  n1908 ) ;
 assign n735 = ( (~ n1938)  &  Ng2912 ) | ( n1938  &  (~ Ng2912) ) ;
 assign Ng24424 = ( n734 ) | ( n735 ) ;
 assign n736 = ( n1858  &  (~ n4869) ) | ( (~ n115)  &  (~ n649)  &  n1858 ) ;
 assign Ng24295 = ( (~ n736) ) ;
 assign n737 = ( n1905  &  Pg3234 ) | ( n1905  &  n1902 ) ;
 assign n738 = ( (~ n1936)  &  Ng3018 ) | ( n1936  &  (~ Ng3018) ) ;
 assign Ng24425 = ( n737 ) | ( n738 ) ;
 assign n739 = ( n1849  &  (~ n4869) ) | ( (~ n118)  &  (~ n654)  &  n1849 ) ;
 assign Ng24336 = ( (~ n739) ) ;
 assign n740 = ( n1840  &  (~ n4869) ) | ( (~ n121)  &  (~ n659)  &  n1840 ) ;
 assign Ng24377 = ( (~ n740) ) ;
 assign n742 = ( (~ Ng2888)  &  n1947 ) | ( Ng2888  &  (~ n1947) ) ;
 assign Ng24423 = ( (~ n714)  &  n742 ) ;
 assign n744 = ( (~ wire1605) ) | ( (~ Ng630) ) ;
 assign n743 = ( wire1605  &  n2706 ) ;
 assign Ng24297 = ( n744  &  Ng738 ) | ( n744  &  n743 ) ;
 assign n745 = ( n1830  &  (~ n4869) ) | ( (~ n124)  &  (~ n662)  &  n1830 ) ;
 assign Ng24418 = ( (~ n745) ) ;
 assign n746 = ( wire1603  &  n2706 ) ;
 assign Ng24298 = ( n707  &  Ng739 ) | ( n707  &  n746 ) ;
 assign n748 = ( (~ wire1605) ) | ( (~ Ng1316) ) ;
 assign n747 = ( wire1605  &  n2705 ) ;
 assign Ng24338 = ( n748  &  Ng1424 ) | ( n748  &  n747 ) ;
 assign n750 = ( (~ wire1605)  &  n3879  &  n3880 ) | ( n3879  &  n3880  &  Ng729 ) ;
 assign n749 = ( (~ wire1603)  &  n383  &  n750 ) | ( n383  &  n750  &  Ng730 ) ;
 assign n752 = ( (~ Ng1315) ) | ( (~ Ng630) ) ;
 assign n751 = ( Ng1315  &  n2706 ) ;
 assign Ng24299 = ( n752  &  Ng737 ) | ( n752  &  n751 ) ;
 assign n753 = ( wire1603  &  n2705 ) ;
 assign Ng24339 = ( n709  &  Ng1425 ) | ( n709  &  n753 ) ;
 assign n755 = ( (~ wire1605) ) | ( (~ Ng2010) ) ;
 assign n754 = ( wire1605  &  n2704 ) ;
 assign Ng24379 = ( n755  &  Ng2118 ) | ( n755  &  n754 ) ;
 assign n757 = ( (~ wire1605)  &  n3876  &  n3877 ) | ( n3876  &  n3877  &  Ng1415 ) ;
 assign n756 = ( (~ wire1603)  &  n433  &  n757 ) | ( n433  &  n757  &  Ng1416 ) ;
 assign n759 = ( (~ Ng1315) ) | ( (~ Ng1316) ) ;
 assign n758 = ( Ng1315  &  n2705 ) ;
 assign Ng24340 = ( n759  &  Ng1423 ) | ( n759  &  n758 ) ;
 assign n760 = ( wire1603  &  n2704 ) ;
 assign Ng24380 = ( n711  &  Ng2119 ) | ( n711  &  n760 ) ;
 assign n762 = ( (~ wire1605) ) | ( (~ Ng2704) ) ;
 assign n761 = ( wire1605  &  n2702 ) ;
 assign Ng24420 = ( n762  &  Ng2812 ) | ( n762  &  n761 ) ;
 assign n764 = ( (~ wire1605)  &  n3873  &  n3874 ) | ( n3873  &  n3874  &  Ng2109 ) ;
 assign n763 = ( (~ wire1603)  &  n478  &  n764 ) | ( n478  &  n764  &  Ng2110 ) ;
 assign n766 = ( (~ Ng1315) ) | ( (~ Ng2010) ) ;
 assign n765 = ( Ng1315  &  n2704 ) ;
 assign Ng24381 = ( n766  &  Ng2117 ) | ( n766  &  n765 ) ;
 assign n767 = ( wire1603  &  n2702 ) ;
 assign Ng24421 = ( n713  &  Ng2813 ) | ( n713  &  n767 ) ;
 assign n769 = ( (~ wire1605)  &  n3870  &  n3871 ) | ( n3870  &  n3871  &  Ng2803 ) ;
 assign n768 = ( (~ wire1603)  &  n513  &  n769 ) | ( n513  &  n769  &  Ng2804 ) ;
 assign n771 = ( (~ Ng1315) ) | ( (~ Ng2704) ) ;
 assign n770 = ( Ng1315  &  n2702 ) ;
 assign Ng24422 = ( n771  &  Ng2811 ) | ( n771  &  n770 ) ;
 assign Ng28313 = ( (~ wire1521)  &  n1527 ) | ( (~ wire1521)  &  Ng3123 ) ;
 assign n772 = ( (~ Ng653)  &  n1945 ) | ( Ng653  &  (~ n1945) ) ;
 assign Ng25140 = ( n772  &  n707 ) ;
 assign n773 = ( (~ Ng1339)  &  n1943 ) | ( Ng1339  &  (~ n1943) ) ;
 assign Ng25151 = ( n773  &  n709 ) ;
 assign n775 = ( (~ n2694)  &  Ng3006 ) | ( n2694  &  (~ Ng3006) ) ;
 assign Ng25177 = ( n775  &  (~ n1905) ) ;
 assign n776 = ( (~ Ng2033)  &  n1941 ) | ( Ng2033  &  (~ n1941) ) ;
 assign Ng25162 = ( n776  &  n711 ) ;
 assign n777 = ( (~ Ng2727)  &  n1939 ) | ( Ng2727  &  (~ n1939) ) ;
 assign Ng25173 = ( n777  &  n713 ) ;
 assign n778 = ( (~ Ng2917)  &  n1937 ) | ( Ng2917  &  (~ n1937) ) ;
 assign Ng25174 = ( (~ n734)  &  n778 ) ;
 assign n780 = ( (~ n1934)  &  Ng2896 ) | ( n1934  &  (~ Ng2896) ) ;
 assign Ng25175 = ( (~ n714)  &  n780 ) ;
 assign n781 = ( (~ Ng3028)  &  n1935 ) | ( Ng3028  &  (~ n1935) ) ;
 assign Ng25176 = ( (~ n737)  &  n781 ) ;
 assign Ng28696 = ( (~ wire1521)  &  n1527 ) | ( (~ wire1521)  &  Ng3125 ) ;
 assign n783 = ( (~ n1927)  &  Ng646 ) | ( n1927  &  (~ Ng646) ) ;
 assign Ng25991 = ( n783  &  n707 ) ;
 assign n784 = ( (~ n1923)  &  Ng1332 ) | ( n1923  &  (~ Ng1332) ) ;
 assign Ng26000 = ( n784  &  n709 ) ;
 assign n785 = ( (~ n1919)  &  Ng2026 ) | ( n1919  &  (~ Ng2026) ) ;
 assign Ng26009 = ( n785  &  n711 ) ;
 assign n786 = ( (~ n1914)  &  Ng2720 ) | ( n1914  &  (~ Ng2720) ) ;
 assign Ng26018 = ( n786  &  n713 ) ;
 assign n787 = ( n1930  &  Ng3002 ) | ( (~ n1930)  &  (~ Ng3002) ) ;
 assign Ng26021 = ( n787  &  (~ n1905) ) ;
 assign n788 = ( (~ n1907)  &  Ng3036 ) | ( n1907  &  (~ Ng3036) ) ;
 assign Ng26022 = ( (~ n737)  &  n788 ) ;
 assign n789 = ( (~ Ng2892)  &  n1933 ) | ( Ng2892  &  (~ n1933) ) ;
 assign Ng26019 = ( (~ n714)  &  n789 ) ;
 assign n790 = ( (~ n1912)  &  Ng2924 ) | ( n1912  &  (~ Ng2924) ) ;
 assign Ng26020 = ( (~ n734)  &  n790 ) ;
 assign n791 = ( n1928  &  Ng88 ) | ( (~ n1928)  &  (~ Ng88) ) ;
 assign n792 = ( n2450 ) | ( n721 ) ;
 assign Ng26678 = ( n791  &  n792 ) ;
 assign n793 = ( n1924  &  Ng776 ) | ( (~ n1924)  &  (~ Ng776) ) ;
 assign Ng26695 = ( n793  &  n792 ) ;
 assign n794 = ( n1920  &  Ng1462 ) | ( (~ n1920)  &  (~ Ng1462) ) ;
 assign Ng26712 = ( n794  &  n792 ) ;
 assign n795 = ( n1915  &  Ng2156 ) | ( (~ n1915)  &  (~ Ng2156) ) ;
 assign Ng26729 = ( n795  &  n792 ) ;
 assign Ng29166 = ( n1620  &  n1621  &  n1622  &  n1623  &  n1624  &  n1625  &  n1626  &  n1627 ) ;
 assign n796 = ( (~ Ng660)  &  n1926 ) | ( Ng660  &  (~ n1926) ) ;
 assign Ng26691 = ( n796  &  n707 ) ;
 assign n797 = ( (~ Ng1346)  &  n1922 ) | ( Ng1346  &  (~ n1922) ) ;
 assign Ng26708 = ( n797  &  n709 ) ;
 assign n798 = ( Ng3013  &  n2695 ) | ( (~ Ng3013)  &  (~ n2695) ) ;
 assign Ng26750 = ( n798  &  (~ n1905) ) ;
 assign n799 = ( (~ Ng2040)  &  n1918 ) | ( Ng2040  &  (~ n1918) ) ;
 assign Ng26725 = ( n799  &  n711 ) ;
 assign n800 = ( (~ Ng2734)  &  n1913 ) | ( Ng2734  &  (~ n1913) ) ;
 assign Ng26742 = ( n800  &  n713 ) ;
 assign n801 = ( (~ Ng2920)  &  n1911 ) | ( Ng2920  &  (~ n1911) ) ;
 assign Ng26746 = ( (~ n734)  &  n801 ) ;
 assign n802 = ( (~ n2699)  &  Ng2903 ) | ( n2699  &  (~ Ng2903) ) ;
 assign Ng26747 = ( (~ n714)  &  n802 ) ;
 assign n803 = ( (~ Ng3032)  &  n1906 ) | ( Ng3032  &  (~ n1906) ) ;
 assign Ng26749 = ( (~ n737)  &  n803 ) ;
 assign n804 = ( (~ n1885)  &  Ng83 ) | ( n1885  &  (~ Ng83) ) ;
 assign Ng27189 = ( n804  &  n792 ) ;
 assign n805 = ( (~ n1881)  &  Ng771 ) | ( n1881  &  (~ Ng771) ) ;
 assign Ng27198 = ( n805  &  n792 ) ;
 assign n806 = ( (~ n1877)  &  Ng1457 ) | ( n1877  &  (~ Ng1457) ) ;
 assign Ng27219 = ( n806  &  n792 ) ;
 assign n807 = ( (~ n1873)  &  Ng2151 ) | ( n1873  &  (~ Ng2151) ) ;
 assign Ng27228 = ( n807  &  n792 ) ;
 assign n808 = ( (~ n1883)  &  Ng672 ) | ( n1883  &  (~ Ng672) ) ;
 assign Ng27197 = ( n808  &  n707 ) ;
 assign n809 = ( (~ n1879)  &  Ng1358 ) | ( n1879  &  (~ Ng1358) ) ;
 assign Ng27218 = ( n809  &  n709 ) ;
 assign n810 = ( (~ n1875)  &  Ng2052 ) | ( n1875  &  (~ Ng2052) ) ;
 assign Ng27227 = ( n810  &  n711 ) ;
 assign n811 = ( (~ n1871)  &  Ng2746 ) | ( n1871  &  (~ Ng2746) ) ;
 assign Ng27236 = ( n811  &  n713 ) ;
 assign n812 = ( n1867  &  Ng3010 ) | ( (~ n1867)  &  (~ Ng3010) ) ;
 assign Ng27239 = ( n812  &  (~ n1905) ) ;
 assign n813 = ( (~ Ng2900)  &  n1869 ) | ( Ng2900  &  (~ n1869) ) ;
 assign Ng27237 = ( (~ n714)  &  n813 ) ;
 assign n814 = ( (~ Ng79)  &  n1884 ) | ( Ng79  &  (~ n1884) ) ;
 assign Ng27683 = ( n814  &  n792 ) ;
 assign n815 = ( (~ Ng767)  &  n1880 ) | ( Ng767  &  (~ n1880) ) ;
 assign Ng27691 = ( n815  &  n792 ) ;
 assign n816 = ( (~ Ng1453)  &  n1876 ) | ( Ng1453  &  (~ n1876) ) ;
 assign Ng27699 = ( n816  &  n792 ) ;
 assign n817 = ( (~ Ng2147)  &  n1872 ) | ( Ng2147  &  (~ n1872) ) ;
 assign Ng27707 = ( n817  &  n792 ) ;
 assign Ng29656 = ( (~ wire1521)  &  n1529  &  Ng185 ) | ( (~ wire1521)  &  n1529  &  n1527 ) ;
 assign n818 = ( (~ Ng666)  &  n1882 ) | ( Ng666  &  (~ n1882) ) ;
 assign Ng27690 = ( n818  &  n707 ) ;
 assign n819 = ( (~ Ng1352)  &  n1878 ) | ( Ng1352  &  (~ n1878) ) ;
 assign Ng27698 = ( n819  &  n709 ) ;
 assign Ng27716 = ( (~ n1905)  &  (~ n2714) ) ;
 assign n821 = ( (~ Ng2046)  &  n1874 ) | ( Ng2046  &  (~ n1874) ) ;
 assign Ng27706 = ( n821  &  n711 ) ;
 assign n822 = ( (~ Ng2740)  &  n1870 ) | ( Ng2740  &  (~ n1870) ) ;
 assign Ng27714 = ( n822  &  n713 ) ;
 assign n823 = ( (~ Ng2908)  &  n1868 ) | ( Ng2908  &  (~ n1868) ) ;
 assign Ng27715 = ( (~ n714)  &  n823 ) ;
 assign n824 = ( (~ n1826)  &  Ng74 ) | ( n1826  &  (~ Ng74) ) ;
 assign Ng28206 = ( n824  &  n792 ) ;
 assign n825 = ( (~ n1816)  &  Ng762 ) | ( n1816  &  (~ Ng762) ) ;
 assign Ng28232 = ( n825  &  n792 ) ;
 assign n826 = ( (~ n1806)  &  Ng1448 ) | ( n1806  &  (~ Ng1448) ) ;
 assign Ng28258 = ( n826  &  n792 ) ;
 assign n827 = ( (~ n1796)  &  Ng2142 ) | ( n1796  &  (~ Ng2142) ) ;
 assign Ng28284 = ( n827  &  n792 ) ;
 assign n828 = ( (~ n2599)  &  Ng679 ) | ( n2599  &  (~ Ng679) ) ;
 assign Ng28231 = ( n828  &  n707 ) ;
 assign n829 = ( (~ n2575)  &  Ng1365 ) | ( n2575  &  (~ Ng1365) ) ;
 assign Ng28257 = ( n829  &  n709 ) ;
 assign n830 = ( (~ n2551)  &  Ng2059 ) | ( n2551  &  (~ Ng2059) ) ;
 assign Ng28283 = ( n830  &  n711 ) ;
 assign n831 = ( (~ n2523)  &  Ng2753 ) | ( n2523  &  (~ Ng2753) ) ;
 assign Ng28309 = ( n831  &  n713 ) ;
 assign n833 = ( n1437  &  n1439  &  n1440 ) ;
 assign n834 = ( n208  &  n1481 ) | ( (~ n208)  &  (~ n1481) ) ;
 assign n832 = ( n833  &  n834 ) ;
 assign n836 = ( n1404  &  n1406  &  n1407 ) ;
 assign n837 = ( n232  &  n1473 ) | ( (~ n232)  &  (~ n1473) ) ;
 assign n835 = ( n836  &  n837 ) ;
 assign n839 = ( n1371  &  n1373  &  n1374 ) ;
 assign n840 = ( n260  &  n1465 ) | ( (~ n260)  &  (~ n1465) ) ;
 assign n838 = ( n839  &  n840 ) ;
 assign n842 = ( n1338  &  n1340  &  n1341 ) ;
 assign n843 = ( n295  &  n1457 ) | ( (~ n295)  &  (~ n1457) ) ;
 assign n841 = ( n842  &  n843 ) ;
 assign n844 = ( (~ Ng70)  &  n1825 ) | ( Ng70  &  (~ n1825) ) ;
 assign Ng28673 = ( n844  &  n792 ) ;
 assign n845 = ( (~ Ng758)  &  n1815 ) | ( Ng758  &  (~ n1815) ) ;
 assign Ng28678 = ( n845  &  n792 ) ;
 assign n846 = ( (~ Ng1444)  &  n1805 ) | ( Ng1444  &  (~ n1805) ) ;
 assign Ng28683 = ( n846  &  n792 ) ;
 assign n847 = ( (~ Ng2138)  &  n1795 ) | ( Ng2138  &  (~ n1795) ) ;
 assign Ng28688 = ( n847  &  n792 ) ;
 assign n848 = ( (~ Ng686)  &  n1734 ) | ( Ng686  &  (~ n1734) ) ;
 assign Ng28677 = ( n848  &  n707 ) ;
 assign n849 = ( (~ Ng1372)  &  n1699 ) | ( Ng1372  &  (~ n1699) ) ;
 assign Ng28682 = ( n849  &  n709 ) ;
 assign n850 = ( (~ Ng2066)  &  n1664 ) | ( Ng2066  &  (~ n1664) ) ;
 assign Ng28687 = ( n850  &  n711 ) ;
 assign n851 = ( (~ Ng2760)  &  n1629 ) | ( Ng2760  &  (~ n1629) ) ;
 assign Ng28692 = ( n851  &  n713 ) ;
 assign n852 = ( (~ n127) ) | ( (~ Ng2257) ) | ( n2680 ) ;
 assign n853 = ( wire1612  &  (~ n1821) ) ;
 assign Ng28674 = ( (~ wire1612)  &  n853 ) | ( n852  &  n853 ) | ( (~ wire1612)  &  Ng448 ) | ( n852  &  Ng448 ) ;
 assign n854 = ( wire1594  &  (~ n1821) ) ;
 assign Ng28675 = ( (~ wire1594)  &  Ng449 ) | ( Ng449  &  n852 ) | ( (~ wire1594)  &  n854 ) | ( n852  &  n854 ) ;
 assign n855 = ( (~ n135) ) | ( (~ Ng2257) ) | ( n2671 ) ;
 assign n856 = ( wire1612  &  (~ n1811) ) ;
 assign Ng28679 = ( (~ wire1612)  &  n856 ) | ( n855  &  n856 ) | ( (~ wire1612)  &  Ng1135 ) | ( n855  &  Ng1135 ) ;
 assign n857 = ( Ng853  &  (~ n1821) ) ;
 assign Ng28676 = ( (~ Ng853)  &  n857 ) | ( n852  &  n857 ) | ( (~ Ng853)  &  Ng447 ) | ( n852  &  Ng447 ) ;
 assign n858 = ( wire1594  &  (~ n1811) ) ;
 assign Ng28680 = ( (~ wire1594)  &  Ng1136 ) | ( Ng1136  &  n855 ) | ( (~ wire1594)  &  n858 ) | ( n855  &  n858 ) ;
 assign n859 = ( (~ n142) ) | ( (~ Ng2257) ) | ( n2662 ) ;
 assign n860 = ( wire1612  &  (~ n1801) ) ;
 assign Ng28684 = ( (~ wire1612)  &  n860 ) | ( n859  &  n860 ) | ( (~ wire1612)  &  Ng1829 ) | ( n859  &  Ng1829 ) ;
 assign n861 = ( Ng853  &  (~ n1811) ) ;
 assign Ng28681 = ( (~ Ng853)  &  n861 ) | ( n855  &  n861 ) | ( (~ Ng853)  &  Ng1134 ) | ( n855  &  Ng1134 ) ;
 assign n862 = ( wire1594  &  (~ n1801) ) ;
 assign Ng28685 = ( (~ wire1594)  &  Ng1830 ) | ( Ng1830  &  n859 ) | ( (~ wire1594)  &  n862 ) | ( n859  &  n862 ) ;
 assign n863 = ( (~ n151) ) | ( (~ Ng2257) ) | ( n2653 ) ;
 assign n864 = ( wire1612  &  (~ n1790) ) ;
 assign Ng28689 = ( (~ wire1612)  &  n864 ) | ( n863  &  n864 ) | ( (~ wire1612)  &  Ng2523 ) | ( n863  &  Ng2523 ) ;
 assign n865 = ( Ng853  &  (~ n1801) ) ;
 assign Ng28686 = ( (~ Ng853)  &  n865 ) | ( n859  &  n865 ) | ( (~ Ng853)  &  Ng1828 ) | ( n859  &  Ng1828 ) ;
 assign n866 = ( wire1594  &  (~ n1790) ) ;
 assign Ng28690 = ( (~ wire1594)  &  Ng2524 ) | ( Ng2524  &  n863 ) | ( (~ wire1594)  &  n866 ) | ( n863  &  n866 ) ;
 assign n867 = ( Ng853  &  (~ n1790) ) ;
 assign Ng28691 = ( (~ Ng853)  &  n867 ) | ( n863  &  n867 ) | ( (~ Ng853)  &  Ng2522 ) | ( n863  &  Ng2522 ) ;
 assign n868 = ( (~ n1619)  &  Ng65 ) | ( n1619  &  (~ Ng65) ) ;
 assign Ng29131 = ( n868  &  n792 ) ;
 assign n869 = ( (~ n1612)  &  Ng753 ) | ( n1612  &  (~ Ng753) ) ;
 assign Ng29139 = ( n869  &  n792 ) ;
 assign n870 = ( (~ n1605)  &  Ng1439 ) | ( n1605  &  (~ Ng1439) ) ;
 assign Ng29147 = ( n870  &  n792 ) ;
 assign n871 = ( (~ n1598)  &  Ng2133 ) | ( n1598  &  (~ Ng2133) ) ;
 assign Ng29155 = ( n871  &  n792 ) ;
 assign n872 = ( (~ Ng692)  &  n1733 ) | ( Ng692  &  (~ n1733) ) ;
 assign Ng29138 = ( n872  &  n707 ) ;
 assign n873 = ( (~ Ng1378)  &  n1698 ) | ( Ng1378  &  (~ n1698) ) ;
 assign Ng29146 = ( n873  &  n709 ) ;
 assign n874 = ( (~ Ng2072)  &  n1663 ) | ( Ng2072  &  (~ n1663) ) ;
 assign Ng29154 = ( n874  &  n711 ) ;
 assign n875 = ( (~ Ng2766)  &  n1628 ) | ( Ng2766  &  (~ n1628) ) ;
 assign Ng29162 = ( n875  &  n713 ) ;
 assign n876 = ( (~ Ng61)  &  n1618 ) | ( Ng61  &  (~ n1618) ) ;
 assign Ng29413 = ( n876  &  n792 ) ;
 assign n877 = ( (~ Ng749)  &  n1611 ) | ( Ng749  &  (~ n1611) ) ;
 assign Ng29420 = ( n877  &  n792 ) ;
 assign n878 = ( (~ Ng1435)  &  n1604 ) | ( Ng1435  &  (~ n1604) ) ;
 assign Ng29427 = ( n878  &  n792 ) ;
 assign n879 = ( (~ Ng2129)  &  n1597 ) | ( Ng2129  &  (~ n1597) ) ;
 assign Ng29446 = ( n879  &  n792 ) ;
 assign n881 = ( (~ wire1612) ) | ( n2495 ) ;
 assign n880 = ( n578  &  (~ n1205)  &  Ng2257 ) ;
 assign Ng29417 = ( n881  &  Ng427 ) | ( n881  &  wire1612  &  n880 ) ;
 assign n882 = ( (~ wire1594) ) | ( n2495 ) ;
 assign Ng29418 = ( n882  &  Ng428 ) | ( n882  &  wire1594  &  n880 ) ;
 assign n884 = ( (~ wire1612) ) | ( n2493 ) ;
 assign n883 = ( n592  &  (~ n1208)  &  Ng2257 ) ;
 assign Ng29424 = ( n884  &  Ng1114 ) | ( n884  &  wire1612  &  n883 ) ;
 assign n885 = ( (~ Ng853) ) | ( n2495 ) ;
 assign Ng29419 = ( n885  &  Ng426 ) | ( n885  &  Ng853  &  n880 ) ;
 assign n886 = ( (~ wire1594) ) | ( n2493 ) ;
 assign Ng29425 = ( n886  &  Ng1115 ) | ( n886  &  wire1594  &  n883 ) ;
 assign n888 = ( (~ wire1612) ) | ( n2491 ) ;
 assign n887 = ( n606  &  (~ n1211)  &  Ng2257 ) ;
 assign Ng29437 = ( n888  &  Ng1808 ) | ( n888  &  wire1612  &  n887 ) ;
 assign n889 = ( (~ Ng853) ) | ( n2493 ) ;
 assign Ng29426 = ( n889  &  Ng1113 ) | ( n889  &  Ng853  &  n883 ) ;
 assign n890 = ( (~ wire1594) ) | ( n2491 ) ;
 assign Ng29438 = ( n890  &  Ng1809 ) | ( n890  &  wire1594  &  n887 ) ;
 assign n892 = ( (~ wire1612) ) | ( n2489 ) ;
 assign n891 = ( n620  &  (~ n1214)  &  Ng2257 ) ;
 assign Ng29450 = ( n892  &  Ng2502 ) | ( n892  &  wire1612  &  n891 ) ;
 assign n893 = ( (~ Ng853) ) | ( n2491 ) ;
 assign Ng29439 = ( n893  &  Ng1807 ) | ( n893  &  Ng853  &  n887 ) ;
 assign n894 = ( (~ wire1594) ) | ( n2489 ) ;
 assign Ng29451 = ( n894  &  Ng2503 ) | ( n894  &  wire1594  &  n891 ) ;
 assign n895 = ( (~ Ng853) ) | ( n2489 ) ;
 assign Ng29452 = ( n895  &  Ng2501 ) | ( n895  &  Ng853  &  n891 ) ;
 assign n896 = ( (~ n1522)  &  Ng56 ) | ( n1522  &  (~ Ng56) ) ;
 assign Ng29627 = ( n896  &  n792 ) ;
 assign n897 = ( (~ n1518)  &  Ng744 ) | ( n1518  &  (~ Ng744) ) ;
 assign Ng29634 = ( n897  &  n792 ) ;
 assign n898 = ( (~ n1514)  &  Ng1430 ) | ( n1514  &  (~ Ng1430) ) ;
 assign Ng29641 = ( n898  &  n792 ) ;
 assign n899 = ( (~ n1510)  &  Ng2124 ) | ( n1510  &  (~ Ng2124) ) ;
 assign Ng29648 = ( n899  &  n792 ) ;
 assign n900 = ( (~ Ng52)  &  n1521 ) | ( Ng52  &  (~ n1521) ) ;
 assign Ng29794 = ( n900  &  n792 ) ;
 assign n901 = ( (~ Ng740)  &  n1517 ) | ( Ng740  &  (~ n1517) ) ;
 assign Ng29798 = ( n901  &  n792 ) ;
 assign n902 = ( (~ Ng1426)  &  n1513 ) | ( Ng1426  &  (~ n1513) ) ;
 assign Ng29802 = ( n902  &  n792 ) ;
 assign n903 = ( (~ Ng2120)  &  n1509 ) | ( Ng2120  &  (~ n1509) ) ;
 assign Ng29806 = ( n903  &  n792 ) ;
 assign n907 = ( n1038 ) | ( n1443 ) ;
 assign n908 = ( n130 ) | ( n1575 ) ;
 assign n904 = ( (~ n542)  &  n907  &  n908 ) | ( n907  &  n908  &  (~ n1038) ) ;
 assign n912 = ( n1042 ) | ( n1410 ) ;
 assign n913 = ( n137 ) | ( n1565 ) ;
 assign n909 = ( (~ n551)  &  n912  &  n913 ) | ( n912  &  n913  &  (~ n1042) ) ;
 assign n917 = ( n1046 ) | ( n1377 ) ;
 assign n918 = ( n144 ) | ( n1555 ) ;
 assign n914 = ( (~ n560)  &  n917  &  n918 ) | ( n917  &  n918  &  (~ n1046) ) ;
 assign n922 = ( n1050 ) | ( n1344 ) ;
 assign n923 = ( n153 ) | ( n1545 ) ;
 assign n919 = ( (~ n567)  &  n922  &  n923 ) | ( n922  &  n923  &  (~ n1050) ) ;
 assign n925 = ( n208  &  n833 ) | ( (~ n208)  &  (~ n833) ) ;
 assign n927 = ( (~ n625)  &  (~ n1448) ) ;
 assign n924 = ( n925  &  n927 ) | ( n925  &  (~ n1264) ) | ( n927  &  (~ n1450) ) | ( (~ n1264)  &  (~ n1450) ) ;
 assign n930 = ( (~ n223)  &  n2117 ) | ( n223  &  (~ n2117) ) ;
 assign n931 = ( Ng101  &  (~ n1448) ) ;
 assign n929 = ( n930  &  n931 ) | ( n930  &  (~ n1264) ) | ( n931  &  (~ n1450) ) | ( (~ n1264)  &  (~ n1450) ) ;
 assign n933 = ( n232  &  n836 ) | ( (~ n232)  &  (~ n836) ) ;
 assign n935 = ( (~ n634)  &  (~ n1415) ) ;
 assign n932 = ( n933  &  n935 ) | ( n933  &  (~ n1267) ) | ( n935  &  (~ n1417) ) | ( (~ n1267)  &  (~ n1417) ) ;
 assign n938 = ( (~ n244)  &  n2116 ) | ( n244  &  (~ n2116) ) ;
 assign n939 = ( Ng109  &  (~ n1448) ) ;
 assign n937 = ( n938  &  n939 ) | ( n938  &  (~ n1264) ) | ( n939  &  (~ n1450) ) | ( (~ n1264)  &  (~ n1450) ) ;
 assign n941 = ( (~ n251)  &  n2084 ) | ( n251  &  (~ n2084) ) ;
 assign n942 = ( Ng789  &  (~ n1415) ) ;
 assign n940 = ( n941  &  n942 ) | ( n941  &  (~ n1267) ) | ( n942  &  (~ n1417) ) | ( (~ n1267)  &  (~ n1417) ) ;
 assign n944 = ( n260  &  n839 ) | ( (~ n260)  &  (~ n839) ) ;
 assign n946 = ( (~ n638)  &  (~ n1382) ) ;
 assign n943 = ( n944  &  n946 ) | ( n944  &  (~ n1270) ) | ( n946  &  (~ n1384) ) | ( (~ n1270)  &  (~ n1384) ) ;
 assign n949 = ( (~ n279)  &  n2083 ) | ( n279  &  (~ n2083) ) ;
 assign n950 = ( Ng797  &  (~ n1415) ) ;
 assign n948 = ( n949  &  n950 ) | ( n949  &  (~ n1267) ) | ( n950  &  (~ n1417) ) | ( (~ n1267)  &  (~ n1417) ) ;
 assign n952 = ( (~ n286)  &  n2051 ) | ( n286  &  (~ n2051) ) ;
 assign n953 = ( Ng1476  &  (~ n1382) ) ;
 assign n951 = ( n952  &  n953 ) | ( n952  &  (~ n1270) ) | ( n953  &  (~ n1384) ) | ( (~ n1270)  &  (~ n1384) ) ;
 assign n955 = ( n295  &  n842 ) | ( (~ n295)  &  (~ n842) ) ;
 assign n957 = ( (~ n642)  &  (~ n1349) ) ;
 assign n954 = ( n955  &  n957 ) | ( n955  &  (~ n1273) ) | ( n957  &  (~ n1351) ) | ( (~ n1273)  &  (~ n1351) ) ;
 assign n960 = ( (~ n321)  &  n2050 ) | ( n321  &  (~ n2050) ) ;
 assign n961 = ( Ng1486  &  (~ n1382) ) ;
 assign n959 = ( n960  &  n961 ) | ( n960  &  (~ n1270) ) | ( n961  &  (~ n1384) ) | ( (~ n1270)  &  (~ n1384) ) ;
 assign n963 = ( (~ n328)  &  n2018 ) | ( n328  &  (~ n2018) ) ;
 assign n964 = ( Ng2170  &  (~ n1349) ) ;
 assign n962 = ( n963  &  n964 ) | ( n963  &  (~ n1273) ) | ( n964  &  (~ n1351) ) | ( (~ n1273)  &  (~ n1351) ) ;
 assign n966 = ( n338  &  n832 ) | ( (~ n338)  &  (~ n832) ) ;
 assign n967 = ( (~ n613)  &  (~ n1448) ) ;
 assign n965 = ( n966  &  n967 ) | ( n966  &  (~ n1264) ) | ( n967  &  (~ n1450) ) | ( (~ n1264)  &  (~ n1450) ) ;
 assign n969 = ( (~ n371)  &  n2017 ) | ( n371  &  (~ n2017) ) ;
 assign n970 = ( Ng2180  &  (~ n1349) ) ;
 assign n968 = ( n969  &  n970 ) | ( n969  &  (~ n1273) ) | ( n970  &  (~ n1351) ) | ( (~ n1273)  &  (~ n1351) ) ;
 assign n972 = ( (~ n376)  &  n2119 ) | ( n376  &  (~ n2119) ) ;
 assign n973 = ( Ng105  &  (~ n1448) ) ;
 assign n971 = ( n972  &  n973 ) | ( n972  &  (~ n1264) ) | ( n973  &  (~ n1450) ) | ( (~ n1264)  &  (~ n1450) ) ;
 assign n975 = ( n388  &  n835 ) | ( (~ n388)  &  (~ n835) ) ;
 assign n976 = ( (~ n627)  &  (~ n1415) ) ;
 assign n974 = ( n975  &  n976 ) | ( n975  &  (~ n1267) ) | ( n976  &  (~ n1417) ) | ( (~ n1267)  &  (~ n1417) ) ;
 assign n978 = ( (~ n426)  &  n2086 ) | ( n426  &  (~ n2086) ) ;
 assign n979 = ( Ng793  &  (~ n1415) ) ;
 assign n977 = ( n978  &  n979 ) | ( n978  &  (~ n1267) ) | ( n979  &  (~ n1417) ) | ( (~ n1267)  &  (~ n1417) ) ;
 assign n981 = ( n438  &  n838 ) | ( (~ n438)  &  (~ n838) ) ;
 assign n982 = ( (~ n636)  &  (~ n1382) ) ;
 assign n980 = ( n981  &  n982 ) | ( n981  &  (~ n1270) ) | ( n982  &  (~ n1384) ) | ( (~ n1270)  &  (~ n1384) ) ;
 assign n984 = ( (~ n471)  &  n2053 ) | ( n471  &  (~ n2053) ) ;
 assign n985 = ( Ng1481  &  (~ n1382) ) ;
 assign n983 = ( n984  &  n985 ) | ( n984  &  (~ n1270) ) | ( n985  &  (~ n1384) ) | ( (~ n1270)  &  (~ n1384) ) ;
 assign n987 = ( n483  &  n841 ) | ( (~ n483)  &  (~ n841) ) ;
 assign n988 = ( (~ n640)  &  (~ n1349) ) ;
 assign n986 = ( n987  &  n988 ) | ( n987  &  (~ n1273) ) | ( n988  &  (~ n1351) ) | ( (~ n1273)  &  (~ n1351) ) ;
 assign n990 = ( (~ n506)  &  n2020 ) | ( n506  &  (~ n2020) ) ;
 assign n991 = ( Ng2175  &  (~ n1349) ) ;
 assign n989 = ( n990  &  n991 ) | ( n990  &  (~ n1273) ) | ( n991  &  (~ n1351) ) | ( (~ n1273)  &  (~ n1351) ) ;
 assign n994 = ( (~ n424) ) | ( n548 ) ;
 assign n993 = ( (~ n548)  &  (~ n1532) ) ;
 assign n992 = ( n424  &  n994  &  (~ n1263) ) | ( n994  &  n993  &  (~ n1263) ) ;
 assign n997 = ( n1532  &  n649 ) ;
 assign n996 = ( n997  &  (~ n1263) ) | ( (~ n1263)  &  (~ n2958) ) ;
 assign n1000 = ( n1532  &  n548 ) ;
 assign n999 = ( n1000  &  (~ n1263) ) | ( (~ n1263)  &  (~ n2959) ) ;
 assign n1004 = ( (~ n381) ) | ( n649 ) ;
 assign n1002 = ( n381  &  n1004  &  (~ n1263) ) | ( n1004  &  (~ n1263)  &  (~ n3738) ) ;
 assign n1005 = ( n997  &  (~ n1263) ) | ( (~ n1263)  &  (~ n2957) ) ;
 assign n1008 = ( (~ n226) ) | ( n548 ) ;
 assign n1007 = ( n226  &  n1008  &  (~ n1263) ) | ( n993  &  n1008  &  (~ n1263) ) ;
 assign n1010 = ( (~ n346) ) | ( n548 ) ;
 assign n1009 = ( n346  &  n1010  &  (~ n1263) ) | ( n993  &  n1010  &  (~ n1263) ) ;
 assign n1012 = ( (~ n462) ) | ( n649 ) ;
 assign n1011 = ( n462  &  n1012  &  (~ n1263) ) | ( n1012  &  (~ n1263)  &  (~ n3738) ) ;
 assign n1015 = ( Pg563 ) | ( n1530 ) | ( Ng559 ) | ( (~ n2727) ) ;
 assign n1013 = ( n1015  &  (~ n1579) ) | ( Ng8284  &  (~ n1262)  &  (~ n1579) ) ;
 assign n1019 = ( (~ n497) ) | ( n654 ) ;
 assign n1017 = ( n497  &  n1019  &  (~ n1260) ) | ( n1019  &  (~ n1260)  &  (~ n3739) ) ;
 assign n1023 = ( (~ n469) ) | ( n557 ) ;
 assign n1022 = ( (~ n557)  &  (~ n1487) ) ;
 assign n1021 = ( n469  &  n1023  &  (~ n1260) ) | ( n1023  &  n1022  &  (~ n1260) ) ;
 assign n1025 = ( n1487  &  n654 ) ;
 assign n1024 = ( n1025  &  (~ n1260) ) | ( (~ n1260)  &  (~ n2939) ) ;
 assign n1028 = ( n1487  &  n557 ) ;
 assign n1027 = ( n1028  &  (~ n1260) ) | ( (~ n1260)  &  (~ n2940) ) ;
 assign n1031 = ( (~ n431) ) | ( n654 ) ;
 assign n1030 = ( n431  &  n1031  &  (~ n1260) ) | ( n1031  &  (~ n1260)  &  (~ n3739) ) ;
 assign n1032 = ( n1025  &  (~ n1260) ) | ( (~ n1260)  &  (~ n2938) ) ;
 assign n1035 = ( (~ n254) ) | ( n557 ) ;
 assign n1034 = ( n254  &  n1035  &  (~ n1260) ) | ( n1022  &  n1035  &  (~ n1260) ) ;
 assign n1037 = ( (~ n396) ) | ( n557 ) ;
 assign n1036 = ( n396  &  n1037  &  (~ n1260) ) | ( n1022  &  n1037  &  (~ n1260) ) ;
 assign n1039 = ( n542  &  (~ n1427) ) | ( (~ n542)  &  n2428 ) | ( (~ n1427)  &  n2428 ) ;
 assign n1038 = ( (~ n534)  &  n538  &  (~ n3988) ) | ( (~ n534)  &  n1039  &  (~ n3988) ) ;
 assign n1043 = ( n551  &  (~ n1394) ) | ( (~ n551)  &  n2393 ) | ( (~ n1394)  &  n2393 ) ;
 assign n1042 = ( (~ n540)  &  n544  &  (~ n3983) ) | ( (~ n540)  &  n1043  &  (~ n3983) ) ;
 assign n1047 = ( n560  &  (~ n1361) ) | ( (~ n560)  &  n2358 ) | ( (~ n1361)  &  n2358 ) ;
 assign n1046 = ( (~ n546)  &  n553  &  (~ n3978) ) | ( (~ n546)  &  n1047  &  (~ n3978) ) ;
 assign n1051 = ( n567  &  (~ n1328) ) | ( (~ n567)  &  n2323 ) | ( (~ n1328)  &  n2323 ) ;
 assign n1050 = ( (~ n555)  &  n562  &  (~ n3973) ) | ( (~ n555)  &  n1051  &  (~ n3973) ) ;
 assign n1056 = ( Pg1249 ) | ( Ng1245 ) | ( (~ n2728) ) ;
 assign n1054 = ( n1056  &  (~ n1494) ) | ( Ng8293  &  (~ n1259)  &  (~ n1494) ) ;
 assign n1059 = ( (~ n542)  &  (~ n1431) ) | ( n1422  &  (~ n1431) ) | ( (~ n1431)  &  (~ n2428) ) ;
 assign n1058 = ( (~ n534)  &  n538  &  (~ n3958) ) | ( (~ n534)  &  n1059  &  (~ n3958) ) ;
 assign n1062 = ( (~ n551)  &  (~ n1398) ) | ( n1389  &  (~ n1398) ) | ( (~ n1398)  &  (~ n2393) ) ;
 assign n1061 = ( (~ n540)  &  n544  &  (~ n3942) ) | ( (~ n540)  &  n1062  &  (~ n3942) ) ;
 assign n1065 = ( (~ n560)  &  (~ n1365) ) | ( n1356  &  (~ n1365) ) | ( (~ n1365)  &  (~ n2358) ) ;
 assign n1064 = ( (~ n546)  &  n553  &  (~ n3926) ) | ( (~ n546)  &  n1065  &  (~ n3926) ) ;
 assign n1068 = ( (~ n567)  &  (~ n1332) ) | ( n1323  &  (~ n1332) ) | ( (~ n1332)  &  (~ n2323) ) ;
 assign n1067 = ( (~ n555)  &  n562  &  (~ n3910) ) | ( (~ n555)  &  n1068  &  (~ n3910) ) ;
 assign n1072 = ( n446  &  n564 ) | ( (~ n446)  &  n3740 ) | ( n564  &  n3740 ) ;
 assign n1070 = ( n1072  &  (~ n1257) ) ;
 assign n1074 = ( n519  &  n659 ) | ( (~ n519)  &  (~ n3741) ) | ( n659  &  (~ n3741) ) ;
 assign n1073 = ( n1074  &  (~ n1257) ) ;
 assign n1076 = ( n504  &  n564 ) | ( (~ n504)  &  n3740 ) | ( n564  &  n3740 ) ;
 assign n1075 = ( n1076  &  (~ n1257) ) ;
 assign n1078 = ( n659  &  (~ n1300) ) ;
 assign n1077 = ( n1078  &  (~ n1257) ) | ( (~ n1257)  &  (~ n2741) ) ;
 assign n1081 = ( n564  &  (~ n1300) ) ;
 assign n1080 = ( n1081  &  (~ n1257) ) | ( (~ n1257)  &  (~ n2742) ) ;
 assign n1084 = ( n476  &  n659 ) | ( (~ n476)  &  (~ n3741) ) | ( n659  &  (~ n3741) ) ;
 assign n1083 = ( n1084  &  (~ n1257) ) ;
 assign n1085 = ( n1078  &  (~ n1257) ) | ( (~ n1257)  &  (~ n2740) ) ;
 assign n1088 = ( n289  &  n564 ) | ( (~ n289)  &  n3740 ) | ( n564  &  n3740 ) ;
 assign n1087 = ( n1088  &  (~ n1257) ) ;
 assign n1091 = ( Pg1943 ) | ( Ng1939 ) | ( (~ n2729) ) ;
 assign n1089 = ( n1091  &  (~ n1311) ) | ( Ng8302  &  (~ n1256)  &  (~ n1311) ) ;
 assign n1094 = ( n1115 ) | ( (~ Ng8311) ) ;
 assign n1093 = ( n1094 ) | ( (~ n3895) ) ;
 assign n1098 = ( n491  &  n569 ) | ( (~ n491)  &  n3742 ) | ( n569  &  n3742 ) ;
 assign n1096 = ( (~ n1094)  &  n1098 ) ;
 assign n1100 = ( n532  &  n662 ) | ( (~ n532)  &  (~ n3743) ) | ( n662  &  (~ n3743) ) ;
 assign n1099 = ( (~ n1094)  &  n1100 ) ;
 assign n1102 = ( n526  &  n569 ) | ( (~ n526)  &  n3742 ) | ( n569  &  n3742 ) ;
 assign n1101 = ( (~ n1094)  &  n1102 ) ;
 assign n1104 = ( n662  &  (~ n1276) ) ;
 assign n1103 = ( (~ n1094)  &  n1104 ) | ( (~ n1094)  &  (~ n2733) ) ;
 assign n1107 = ( n569  &  (~ n1276) ) ;
 assign n1106 = ( (~ n1094)  &  n1107 ) | ( (~ n1094)  &  (~ n2734) ) ;
 assign n1110 = ( n511  &  n662 ) | ( (~ n511)  &  (~ n3743) ) | ( n662  &  (~ n3743) ) ;
 assign n1109 = ( (~ n1094)  &  n1110 ) ;
 assign n1111 = ( (~ n1094)  &  n1104 ) | ( (~ n1094)  &  (~ n2732) ) ;
 assign n1115 = ( Pg2637 ) | ( Ng2633 ) | ( (~ n2730) ) ;
 assign n1113 = ( n1115  &  (~ n1287) ) | ( Ng8311  &  (~ n1254)  &  (~ n1287) ) ;
 assign n1118 = ( Ng2874  &  Ng2981 ) | ( (~ Ng2874)  &  (~ Ng2981) ) ;
 assign n1119 = ( Ng2978  &  Ng2975 ) | ( (~ Ng2978)  &  (~ Ng2975) ) ;
 assign n1120 = ( (~ Ng2874)  &  Ng2981 ) | ( Ng2874  &  (~ Ng2981) ) ;
 assign n1121 = ( (~ Ng2978)  &  Ng2975 ) | ( Ng2978  &  (~ Ng2975) ) ;
 assign n1117 = ( n1118  &  n1120 ) | ( n1119  &  n1120 ) | ( n1118  &  n1121 ) | ( n1119  &  n1121 ) ;
 assign n1123 = ( Ng2972  &  Ng2969 ) | ( (~ Ng2972)  &  (~ Ng2969) ) ;
 assign n1124 = ( Ng2966  &  Ng2963 ) | ( (~ Ng2966)  &  (~ Ng2963) ) ;
 assign n1125 = ( (~ Ng2972)  &  Ng2969 ) | ( Ng2972  &  (~ Ng2969) ) ;
 assign n1126 = ( (~ Ng2966)  &  Ng2963 ) | ( Ng2966  &  (~ Ng2963) ) ;
 assign n1122 = ( n1123  &  n1125 ) | ( n1124  &  n1125 ) | ( n1123  &  n1126 ) | ( n1124  &  n1126 ) ;
 assign n1128 = ( Ng2959  &  Ng2956 ) | ( (~ Ng2959)  &  (~ Ng2956) ) ;
 assign n1129 = ( Ng2953  &  Ng2947 ) | ( (~ Ng2953)  &  (~ Ng2947) ) ;
 assign n1130 = ( (~ Ng2959)  &  Ng2956 ) | ( Ng2959  &  (~ Ng2956) ) ;
 assign n1131 = ( (~ Ng2953)  &  Ng2947 ) | ( Ng2953  &  (~ Ng2947) ) ;
 assign n1127 = ( n1128  &  n1130 ) | ( n1129  &  n1130 ) | ( n1128  &  n1131 ) | ( n1129  &  n1131 ) ;
 assign n1133 = ( Ng2944  &  Ng2941 ) | ( (~ Ng2944)  &  (~ Ng2941) ) ;
 assign n1134 = ( Ng2938  &  Ng2935 ) | ( (~ Ng2938)  &  (~ Ng2935) ) ;
 assign n1135 = ( (~ Ng2944)  &  Ng2941 ) | ( Ng2944  &  (~ Ng2941) ) ;
 assign n1136 = ( (~ Ng2938)  &  Ng2935 ) | ( Ng2938  &  (~ Ng2935) ) ;
 assign n1132 = ( n1133  &  n1135 ) | ( n1134  &  n1135 ) | ( n1133  &  n1136 ) | ( n1134  &  n1136 ) ;
 assign n1149 = ( n1000  &  (~ n1263) ) | ( (~ n1263)  &  (~ n2955) ) ;
 assign n1151 = ( n997  &  (~ n1263) ) | ( (~ n1263)  &  (~ n2956) ) ;
 assign n1154 = ( n992  &  n1011 ) | ( (~ n992)  &  (~ n1011) ) ;
 assign n1155 = ( n1002  &  n1009 ) | ( (~ n1002)  &  (~ n1009) ) ;
 assign n1156 = ( (~ n992)  &  n1011 ) | ( n992  &  (~ n1011) ) ;
 assign n1157 = ( (~ n1002)  &  n1009 ) | ( n1002  &  (~ n1009) ) ;
 assign n1153 = ( n1154  &  n1156 ) | ( n1155  &  n1156 ) | ( n1154  &  n1157 ) | ( n1155  &  n1157 ) ;
 assign n1159 = ( n1005  &  n1007 ) | ( (~ n1005)  &  (~ n1007) ) ;
 assign n1160 = ( n996  &  n999 ) | ( (~ n996)  &  (~ n999) ) ;
 assign n1161 = ( (~ n1005)  &  n1007 ) | ( n1005  &  (~ n1007) ) ;
 assign n1162 = ( (~ n996)  &  n999 ) | ( n996  &  (~ n999) ) ;
 assign n1158 = ( n1159  &  n1161 ) | ( n1160  &  n1161 ) | ( n1159  &  n1162 ) | ( n1160  &  n1162 ) ;
 assign n1163 = ( n1028  &  (~ n1260) ) | ( (~ n1260)  &  (~ n2936) ) ;
 assign n1165 = ( n1025  &  (~ n1260) ) | ( (~ n1260)  &  (~ n2937) ) ;
 assign n1168 = ( n1030  &  n1036 ) | ( (~ n1030)  &  (~ n1036) ) ;
 assign n1169 = ( n1017  &  n1021 ) | ( (~ n1017)  &  (~ n1021) ) ;
 assign n1170 = ( (~ n1030)  &  n1036 ) | ( n1030  &  (~ n1036) ) ;
 assign n1171 = ( (~ n1017)  &  n1021 ) | ( n1017  &  (~ n1021) ) ;
 assign n1167 = ( n1168  &  n1170 ) | ( n1169  &  n1170 ) | ( n1168  &  n1171 ) | ( n1169  &  n1171 ) ;
 assign n1173 = ( n1032  &  n1034 ) | ( (~ n1032)  &  (~ n1034) ) ;
 assign n1174 = ( n1024  &  n1027 ) | ( (~ n1024)  &  (~ n1027) ) ;
 assign n1175 = ( (~ n1032)  &  n1034 ) | ( n1032  &  (~ n1034) ) ;
 assign n1176 = ( (~ n1024)  &  n1027 ) | ( n1024  &  (~ n1027) ) ;
 assign n1172 = ( n1173  &  n1175 ) | ( n1174  &  n1175 ) | ( n1173  &  n1176 ) | ( n1174  &  n1176 ) ;
 assign n1177 = ( n1081  &  (~ n1257) ) | ( (~ n1257)  &  (~ n2738) ) ;
 assign n1179 = ( n1078  &  (~ n1257) ) | ( (~ n1257)  &  (~ n2739) ) ;
 assign n1182 = ( n1070  &  n1083 ) | ( (~ n1070)  &  (~ n1083) ) ;
 assign n1183 = ( n1073  &  n1075 ) | ( (~ n1073)  &  (~ n1075) ) ;
 assign n1184 = ( (~ n1070)  &  n1083 ) | ( n1070  &  (~ n1083) ) ;
 assign n1185 = ( (~ n1073)  &  n1075 ) | ( n1073  &  (~ n1075) ) ;
 assign n1181 = ( n1182  &  n1184 ) | ( n1183  &  n1184 ) | ( n1182  &  n1185 ) | ( n1183  &  n1185 ) ;
 assign n1187 = ( n1085  &  n1087 ) | ( (~ n1085)  &  (~ n1087) ) ;
 assign n1188 = ( n1077  &  n1080 ) | ( (~ n1077)  &  (~ n1080) ) ;
 assign n1189 = ( (~ n1085)  &  n1087 ) | ( n1085  &  (~ n1087) ) ;
 assign n1190 = ( (~ n1077)  &  n1080 ) | ( n1077  &  (~ n1080) ) ;
 assign n1186 = ( n1187  &  n1189 ) | ( n1188  &  n1189 ) | ( n1187  &  n1190 ) | ( n1188  &  n1190 ) ;
 assign n1191 = ( (~ n1094)  &  n1107 ) | ( (~ n1094)  &  (~ n2726) ) ;
 assign n1193 = ( (~ n1094)  &  n1104 ) | ( (~ n1094)  &  (~ n2731) ) ;
 assign n1196 = ( n1096  &  n1109 ) | ( (~ n1096)  &  (~ n1109) ) ;
 assign n1197 = ( n1099  &  n1101 ) | ( (~ n1099)  &  (~ n1101) ) ;
 assign n1198 = ( (~ n1096)  &  n1109 ) | ( n1096  &  (~ n1109) ) ;
 assign n1199 = ( (~ n1099)  &  n1101 ) | ( n1099  &  (~ n1101) ) ;
 assign n1195 = ( n1196  &  n1198 ) | ( n1197  &  n1198 ) | ( n1196  &  n1199 ) | ( n1197  &  n1199 ) ;
 assign n1201 = ( (~ n1111)  &  n1093 ) | ( n1111  &  (~ n1093) ) ;
 assign n1202 = ( n1103  &  n1106 ) | ( (~ n1103)  &  (~ n1106) ) ;
 assign n1203 = ( n1093  &  n1111 ) | ( (~ n1093)  &  (~ n1111) ) ;
 assign n1204 = ( (~ n1103)  &  n1106 ) | ( n1103  &  (~ n1106) ) ;
 assign n1200 = ( n1201  &  n1203 ) | ( n1202  &  n1203 ) | ( n1201  &  n1204 ) | ( n1202  &  n1204 ) ;
 assign n1207 = ( (~ n587) ) | ( (~ n1206) ) | ( n2429 ) ;
 assign n1206 = ( (~ n613)  &  (~ n625)  &  n1820 ) ;
 assign n1205 = ( n1207  &  n1206 ) | ( n1207  &  n587 ) ;
 assign n1210 = ( (~ n601) ) | ( (~ n1209) ) | ( n2394 ) ;
 assign n1209 = ( (~ n627)  &  (~ n634)  &  n1810 ) ;
 assign n1208 = ( n1210  &  n1209 ) | ( n1210  &  n601 ) ;
 assign n1213 = ( (~ n615) ) | ( (~ n1212) ) | ( n2359 ) ;
 assign n1212 = ( (~ n636)  &  (~ n638)  &  n1800 ) ;
 assign n1211 = ( n1213  &  n1212 ) | ( n1213  &  n615 ) ;
 assign n1216 = ( (~ n629) ) | ( (~ n1215) ) | ( n2324 ) ;
 assign n1215 = ( (~ n640)  &  (~ n642)  &  n1789 ) ;
 assign n1214 = ( n1216  &  n1215 ) | ( n1216  &  n629 ) ;
 assign Ng19048 = ( (~ n629) ) ;
 assign Ng19036 = ( (~ n615) ) ;
 assign Ng19024 = ( (~ n601) ) ;
 assign Ng19012 = ( (~ n587) ) ;
 assign n1217 = ( (~ Ng2584)  &  n1284 ) | ( n1284  &  n1283 ) ;
 assign Ng30989 = ( (~ n1217) ) ;
 assign n1218 = ( (~ n677)  &  n1191 ) | ( (~ n677)  &  n1287 ) | ( n1191  &  (~ n3748) ) | ( n1287  &  (~ n3748) ) ;
 assign Ng30987 = ( (~ n1218) ) ;
 assign n1219 = ( (~ n677)  &  n1193 ) | ( (~ n677)  &  n1287 ) | ( n1193  &  (~ n3749) ) | ( n1287  &  (~ n3749) ) ;
 assign Ng30986 = ( (~ n1219) ) ;
 assign n1220 = ( (~ n677)  &  n1290 ) | ( n1290  &  (~ n3750) ) ;
 assign Ng30985 = ( (~ n1220) ) ;
 assign n1221 = ( (~ n677)  &  n1290 ) | ( n1290  &  (~ n3751) ) ;
 assign Ng30984 = ( (~ n1221) ) ;
 assign n1222 = ( (~ n677)  &  (~ n1253) ) | ( (~ n1253)  &  (~ n3752) ) ;
 assign Ng30983 = ( (~ n1222) ) ;
 assign n1223 = ( (~ n677)  &  (~ n1113) ) | ( (~ n1113)  &  (~ n3754) ) ;
 assign Ng30982 = ( (~ n1223) ) ;
 assign n1224 = ( (~ n677)  &  (~ n1113) ) | ( (~ n1113)  &  (~ n3755) ) ;
 assign Ng30981 = ( (~ n1224) ) ;
 assign n1225 = ( (~ n677)  &  (~ n1253) ) | ( (~ n1253)  &  (~ n3756) ) ;
 assign Ng30980 = ( (~ n1225) ) ;
 assign n1226 = ( (~ Ng1890)  &  n1308 ) | ( n1308  &  n1307 ) ;
 assign Ng30940 = ( (~ n1226) ) ;
 assign n1227 = ( (~ n673)  &  n1177 ) | ( (~ n673)  &  n1311 ) | ( n1177  &  (~ n3762) ) | ( n1311  &  (~ n3762) ) ;
 assign Ng30915 = ( (~ n1227) ) ;
 assign n1228 = ( (~ n673)  &  n1179 ) | ( (~ n673)  &  n1311 ) | ( n1179  &  (~ n3763) ) | ( n1311  &  (~ n3763) ) ;
 assign Ng30914 = ( (~ n1228) ) ;
 assign n1229 = ( (~ n673)  &  n1314 ) | ( n1314  &  (~ n3764) ) ;
 assign Ng30913 = ( (~ n1229) ) ;
 assign n1230 = ( (~ n673)  &  n1314 ) | ( n1314  &  (~ n3765) ) ;
 assign Ng30912 = ( (~ n1230) ) ;
 assign n1231 = ( (~ n673)  &  (~ n1255) ) | ( (~ n1255)  &  (~ n3766) ) ;
 assign Ng30911 = ( (~ n1231) ) ;
 assign n1232 = ( (~ n673)  &  (~ n1089) ) | ( (~ n1089)  &  (~ n3768) ) ;
 assign Ng30910 = ( (~ n1232) ) ;
 assign n1233 = ( (~ n673)  &  (~ n1089) ) | ( (~ n1089)  &  (~ n3769) ) ;
 assign Ng30909 = ( (~ n1233) ) ;
 assign n1234 = ( (~ n673)  &  (~ n1255) ) | ( (~ n1255)  &  (~ n3770) ) ;
 assign Ng30908 = ( (~ n1234) ) ;
 assign n1235 = ( (~ Ng1196)  &  n1491 ) | ( n1491  &  n1490 ) ;
 assign Ng30119 = ( (~ n1235) ) ;
 assign n1236 = ( (~ n669)  &  n1163 ) | ( (~ n669)  &  n1494 ) | ( n1163  &  (~ n3828) ) | ( n1494  &  (~ n3828) ) ;
 assign Ng29979 = ( (~ n1236) ) ;
 assign n1237 = ( (~ n669)  &  n1165 ) | ( (~ n669)  &  n1494 ) | ( n1165  &  (~ n3829) ) | ( n1494  &  (~ n3829) ) ;
 assign Ng29978 = ( (~ n1237) ) ;
 assign n1238 = ( (~ n669)  &  n1497 ) | ( n1497  &  (~ n3830) ) ;
 assign Ng29977 = ( (~ n1238) ) ;
 assign n1239 = ( (~ n669)  &  n1497 ) | ( n1497  &  (~ n3831) ) ;
 assign Ng29976 = ( (~ n1239) ) ;
 assign n1240 = ( (~ n669)  &  (~ n1258) ) | ( (~ n1258)  &  (~ n3832) ) ;
 assign Ng29975 = ( (~ n1240) ) ;
 assign n1241 = ( (~ n669)  &  (~ n1054) ) | ( (~ n1054)  &  (~ n3833) ) ;
 assign Ng29974 = ( (~ n1241) ) ;
 assign n1242 = ( (~ n669)  &  (~ n1054) ) | ( (~ n1054)  &  (~ n3834) ) ;
 assign Ng29973 = ( (~ n1242) ) ;
 assign n1243 = ( (~ n669)  &  (~ n1258) ) | ( (~ n1258)  &  (~ n3835) ) ;
 assign Ng29972 = ( (~ n1243) ) ;
 assign n1244 = ( (~ Ng510)  &  n1536 ) | ( n1536  &  n1535 ) ;
 assign Ng29655 = ( (~ n1244) ) ;
 assign n1245 = ( (~ n665)  &  n1149 ) | ( (~ n665)  &  n1579 ) | ( n1149  &  (~ n3840) ) | ( n1579  &  (~ n3840) ) ;
 assign Ng29460 = ( (~ n1245) ) ;
 assign n1246 = ( (~ n665)  &  n1151 ) | ( (~ n665)  &  n1579 ) | ( n1151  &  (~ n3841) ) | ( n1579  &  (~ n3841) ) ;
 assign Ng29459 = ( (~ n1246) ) ;
 assign n1247 = ( (~ n665)  &  n1582 ) | ( n1582  &  (~ n3842) ) ;
 assign Ng29458 = ( (~ n1247) ) ;
 assign n1248 = ( (~ n665)  &  n1582 ) | ( n1582  &  (~ n3843) ) ;
 assign Ng29457 = ( (~ n1248) ) ;
 assign n1249 = ( (~ n665)  &  (~ n1261) ) | ( (~ n1261)  &  (~ n3844) ) ;
 assign Ng29456 = ( (~ n1249) ) ;
 assign n1250 = ( (~ n665)  &  (~ n1013) ) | ( (~ n1013)  &  (~ n3845) ) ;
 assign Ng29455 = ( (~ n1250) ) ;
 assign n1251 = ( (~ n665)  &  (~ n1013) ) | ( (~ n1013)  &  (~ n3846) ) ;
 assign Ng29454 = ( (~ n1251) ) ;
 assign n1252 = ( (~ n665)  &  (~ n1261) ) | ( (~ n1261)  &  (~ n3847) ) ;
 assign Ng29453 = ( (~ n1252) ) ;
 assign Ng13466 = ( (~ Ng2366) ) ;
 assign Ng13465 = ( (~ Ng2364) ) ;
 assign Ng13464 = ( (~ Ng2362) ) ;
 assign Ng13463 = ( (~ Ng2360) ) ;
 assign Ng13462 = ( (~ Ng2358) ) ;
 assign Ng13461 = ( (~ Ng2356) ) ;
 assign Ng13460 = ( (~ Ng2354) ) ;
 assign Ng13459 = ( (~ Ng2528) ) ;
 assign Ng13458 = ( (~ Ng2526) ) ;
 assign Ng11576 = ( (~ Ng2165) ) ;
 assign Ng11575 = ( (~ Ng2170) ) ;
 assign Ng11574 = ( (~ Ng2175) ) ;
 assign Ng11573 = ( (~ Ng2180) ) ;
 assign Ng11572 = ( (~ Ng2185) ) ;
 assign Ng11592 = ( (~ Ng2190) ) ;
 assign Ng11591 = ( (~ Ng2195) ) ;
 assign Ng11590 = ( (~ Ng2200) ) ;
 assign Ng13450 = ( (~ Ng1672) ) ;
 assign Ng13449 = ( (~ Ng1670) ) ;
 assign Ng13448 = ( (~ Ng1668) ) ;
 assign Ng13447 = ( (~ Ng1666) ) ;
 assign Ng13446 = ( (~ Ng1664) ) ;
 assign Ng13445 = ( (~ Ng1662) ) ;
 assign Ng13444 = ( (~ Ng1660) ) ;
 assign Ng13443 = ( (~ Ng1834) ) ;
 assign Ng13442 = ( (~ Ng1832) ) ;
 assign Ng11549 = ( (~ Ng1471) ) ;
 assign Ng11548 = ( (~ Ng1476) ) ;
 assign Ng11547 = ( (~ Ng1481) ) ;
 assign Ng11546 = ( (~ Ng1486) ) ;
 assign Ng11545 = ( (~ Ng1491) ) ;
 assign Ng11565 = ( (~ Ng1496) ) ;
 assign Ng11564 = ( (~ Ng1501) ) ;
 assign Ng11563 = ( (~ Ng1506) ) ;
 assign Ng13434 = ( (~ Ng978) ) ;
 assign Ng13433 = ( (~ Ng976) ) ;
 assign Ng13432 = ( (~ Ng974) ) ;
 assign Ng13431 = ( (~ Ng972) ) ;
 assign Ng13430 = ( (~ Ng970) ) ;
 assign Ng13429 = ( (~ Ng968) ) ;
 assign Ng13428 = ( (~ Ng966) ) ;
 assign Ng13427 = ( (~ Ng1140) ) ;
 assign Ng13426 = ( (~ Ng1138) ) ;
 assign Ng11522 = ( (~ Ng785) ) ;
 assign Ng11521 = ( (~ Ng789) ) ;
 assign Ng11520 = ( (~ Ng793) ) ;
 assign Ng11519 = ( (~ Ng797) ) ;
 assign Ng11518 = ( (~ Ng801) ) ;
 assign Ng11538 = ( (~ Ng805) ) ;
 assign Ng11537 = ( (~ Ng809) ) ;
 assign Ng11536 = ( (~ Ng813) ) ;
 assign Ng13418 = ( (~ Ng291) ) ;
 assign Ng13417 = ( (~ Ng289) ) ;
 assign Ng13416 = ( (~ Ng287) ) ;
 assign Ng13415 = ( (~ Ng285) ) ;
 assign Ng13414 = ( (~ Ng283) ) ;
 assign Ng13413 = ( (~ Ng281) ) ;
 assign Ng13412 = ( (~ Ng279) ) ;
 assign Ng13411 = ( (~ Ng453) ) ;
 assign Ng13410 = ( (~ Ng451) ) ;
 assign Ng11495 = ( (~ Ng97) ) ;
 assign Ng11494 = ( (~ Ng101) ) ;
 assign Ng11493 = ( (~ Ng105) ) ;
 assign Ng11492 = ( (~ Ng109) ) ;
 assign Ng11491 = ( (~ Ng113) ) ;
 assign Ng11511 = ( (~ Ng117) ) ;
 assign Ng11510 = ( (~ Ng121) ) ;
 assign Ng11509 = ( (~ Ng125) ) ;
 assign n1254 = ( (~ wire1605)  &  n1276  &  n1293 ) | ( n1276  &  n1293  &  Ng2809 ) ;
 assign n1253 = ( n1094  &  (~ n1287) ) | ( n1254  &  (~ n1287) ) ;
 assign n1256 = ( (~ wire1605)  &  n1300  &  n1316 ) | ( n1300  &  n1316  &  Ng2115 ) ;
 assign n1257 = ( n1091 ) | ( (~ Ng8302) ) ;
 assign n1255 = ( n1256  &  (~ n1311) ) | ( n1257  &  (~ n1311) ) ;
 assign n1259 = ( (~ wire1605)  &  (~ n1487)  &  n1500 ) | ( (~ n1487)  &  n1500  &  Ng1421 ) ;
 assign n1260 = ( n1056 ) | ( (~ Ng8293) ) ;
 assign n1258 = ( n1259  &  (~ n1494) ) | ( n1260  &  (~ n1494) ) ;
 assign n1262 = ( (~ wire1605)  &  (~ n1532)  &  n1585 ) | ( (~ n1532)  &  n1585  &  Ng735 ) ;
 assign n1263 = ( n1015 ) | ( (~ Ng8284) ) ;
 assign n1261 = ( n1262  &  (~ n1579) ) | ( n1263  &  (~ n1579) ) ;
 assign n1264 = ( (~ n1448)  &  (~ n1450) ) | ( (~ n1450)  &  (~ n1481) ) ;
 assign n1267 = ( (~ n1415)  &  (~ n1417) ) | ( (~ n1417)  &  (~ n1473) ) ;
 assign n1270 = ( (~ n1382)  &  (~ n1384) ) | ( (~ n1384)  &  (~ n1465) ) ;
 assign n1273 = ( (~ n1349)  &  (~ n1351) ) | ( (~ n1351)  &  (~ n1457) ) ;
 assign n1282 = ( n513 ) | ( n458 ) | ( n536 ) | ( n374 ) | ( n333 ) | ( n417 ) ;
 assign n1276 = ( (~ n331) ) | ( (~ n491) ) | ( (~ n511) ) | ( (~ n526) ) | ( n1282 ) | ( (~ n3746) ) ;
 assign n1284 = ( (~ Ng2631)  &  n3900 ) | ( n3898  &  n3900 ) ;
 assign n1283 = ( n1195  &  n1200 ) | ( (~ n1195)  &  (~ n1200) ) ;
 assign n1287 = ( n677 ) | ( (~ n679) ) ;
 assign n1290 = ( (~ n1115) ) | ( n1287 ) ;
 assign n1293 = ( (~ wire1603)  &  (~ Ng1315) ) | ( (~ Ng1315)  &  Ng2810 ) | ( (~ wire1603)  &  Ng2808 ) | ( Ng2810  &  Ng2808 ) ;
 assign n1306 = ( n478 ) | ( n408 ) | ( n528 ) | ( n324 ) | ( n291 ) | ( n367 ) ;
 assign n1300 = ( (~ n289) ) | ( (~ n446) ) | ( (~ n476) ) | ( (~ n504) ) | ( n1306 ) | ( (~ n3760) ) ;
 assign n1308 = ( (~ Ng1937)  &  n3907 ) | ( n3905  &  n3907 ) ;
 assign n1307 = ( n1181  &  n1186 ) | ( (~ n1181)  &  (~ n1186) ) ;
 assign n1311 = ( n673 ) | ( (~ n675) ) ;
 assign n1314 = ( (~ n1091) ) | ( n1311 ) ;
 assign n1316 = ( (~ wire1603)  &  (~ Ng1315) ) | ( (~ Ng1315)  &  Ng2116 ) | ( (~ wire1603)  &  Ng2114 ) | ( Ng2116  &  Ng2114 ) ;
 assign n1324 = ( n2003  &  n2006 ) | ( (~ n2005)  &  n2006 ) | ( n2003  &  n2008 ) | ( (~ n2005)  &  n2008 ) ;
 assign n1325 = ( n414  &  Ng2190 ) | ( (~ n414)  &  (~ Ng2190) ) ;
 assign n1323 = ( (~ n1329)  &  (~ n3783) ) | ( n1324  &  n1325  &  (~ n1329) ) ;
 assign n1329 = ( n530 ) | ( (~ Ng2257) ) ;
 assign n1330 = ( n1325 ) | ( n1334 ) | ( n2002 ) | ( n2003 ) | ( (~ n2005) ) | ( n2006 ) | ( n2008 ) | ( n2319 ) ;
 assign n1328 = ( n1329  &  (~ n2324) ) | ( n1330  &  (~ n2324) ) ;
 assign n1333 = ( n1996  &  n2000 ) | ( n1998  &  n2000 ) | ( n1996  &  n2002 ) | ( n1998  &  n2002 ) ;
 assign n1334 = ( (~ n295)  &  n642 ) | ( n295  &  (~ n642) ) ;
 assign n1332 = ( (~ n1329)  &  (~ n3776) ) | ( (~ n1329)  &  n1333  &  n1334 ) ;
 assign n1339 = ( n2009  &  (~ n2020)  &  (~ n2327) ) ;
 assign n1338 = ( n414  &  n1339 ) | ( n1339  &  (~ n1457) ) ;
 assign n1340 = ( n265  &  n1457 ) | ( (~ n265)  &  (~ n1457) ) ;
 assign n1341 = ( (~ n414)  &  (~ n450) ) | ( (~ n414)  &  n1457 ) | ( n450  &  n1457 ) ;
 assign n1343 = ( (~ n1545)  &  (~ n2320) ) ;
 assign n1344 = ( (~ n555)  &  n567 ) ;
 assign n1342 = ( n562  &  n1343  &  n1344 ) ;
 assign n1345 = ( (~ n177)  &  n1342 ) | ( (~ n177)  &  (~ n1545)  &  (~ n1546) ) ;
 assign n1349 = ( n555  &  n923  &  (~ n1345) ) | ( n923  &  (~ n1345)  &  (~ n2324) ) ;
 assign n1352 = ( n1889  &  n1457 ) ;
 assign n1351 = ( n1349  &  n1352 ) | ( n1349  &  (~ n2747) ) ;
 assign n1357 = ( n2036  &  n2039 ) | ( (~ n2038)  &  n2039 ) | ( n2036  &  n2041 ) | ( (~ n2038)  &  n2041 ) ;
 assign n1358 = ( n364  &  Ng1496 ) | ( (~ n364)  &  (~ Ng1496) ) ;
 assign n1356 = ( (~ n1362)  &  (~ n3796) ) | ( n1357  &  n1358  &  (~ n1362) ) ;
 assign n1362 = ( n517 ) | ( (~ Ng2257) ) ;
 assign n1363 = ( n1358 ) | ( n1367 ) | ( n2035 ) | ( n2036 ) | ( (~ n2038) ) | ( n2039 ) | ( n2041 ) | ( n2354 ) ;
 assign n1361 = ( n1362  &  (~ n2359) ) | ( n1363  &  (~ n2359) ) ;
 assign n1366 = ( n2029  &  n2033 ) | ( n2031  &  n2033 ) | ( n2029  &  n2035 ) | ( n2031  &  n2035 ) ;
 assign n1367 = ( (~ n260)  &  n638 ) | ( n260  &  (~ n638) ) ;
 assign n1365 = ( (~ n1362)  &  (~ n3789) ) | ( (~ n1362)  &  n1366  &  n1367 ) ;
 assign n1372 = ( n2042  &  (~ n2053)  &  (~ n2362) ) ;
 assign n1371 = ( n364  &  n1372 ) | ( n1372  &  (~ n1465) ) ;
 assign n1373 = ( n237  &  n1465 ) | ( (~ n237)  &  (~ n1465) ) ;
 assign n1374 = ( (~ n364)  &  (~ n400) ) | ( (~ n364)  &  n1465 ) | ( n400  &  n1465 ) ;
 assign n1376 = ( (~ n1555)  &  (~ n2355) ) ;
 assign n1377 = ( (~ n546)  &  n560 ) ;
 assign n1375 = ( n553  &  n1376  &  n1377 ) ;
 assign n1378 = ( (~ n173)  &  n1375 ) | ( (~ n173)  &  (~ n1555)  &  (~ n1556) ) ;
 assign n1382 = ( n546  &  n918  &  (~ n1378) ) | ( n918  &  (~ n1378)  &  (~ n2359) ) ;
 assign n1385 = ( n1893  &  n1465 ) ;
 assign n1384 = ( n1382  &  n1385 ) | ( n1382  &  (~ n2767) ) ;
 assign n1390 = ( n2069  &  n2072 ) | ( (~ n2071)  &  n2072 ) | ( n2069  &  n2074 ) | ( (~ n2071)  &  n2074 ) ;
 assign n1391 = ( n314  &  Ng805 ) | ( (~ n314)  &  (~ Ng805) ) ;
 assign n1389 = ( (~ n1395)  &  (~ n3809) ) | ( n1390  &  n1391  &  (~ n1395) ) ;
 assign n1395 = ( n495 ) | ( (~ Ng2257) ) ;
 assign n1396 = ( n1391 ) | ( n1400 ) | ( n2068 ) | ( n2069 ) | ( (~ n2071) ) | ( n2072 ) | ( n2074 ) | ( n2389 ) ;
 assign n1394 = ( n1395  &  (~ n2394) ) | ( n1396  &  (~ n2394) ) ;
 assign n1399 = ( n2062  &  n2066 ) | ( n2064  &  n2066 ) | ( n2062  &  n2068 ) | ( n2064  &  n2068 ) ;
 assign n1400 = ( (~ n232)  &  n634 ) | ( n232  &  (~ n634) ) ;
 assign n1398 = ( (~ n1395)  &  (~ n3802) ) | ( (~ n1395)  &  n1399  &  n1400 ) ;
 assign n1405 = ( n2075  &  (~ n2086)  &  (~ n2397) ) ;
 assign n1404 = ( n314  &  n1405 ) | ( n1405  &  (~ n1473) ) ;
 assign n1406 = ( n214  &  n1473 ) | ( (~ n214)  &  (~ n1473) ) ;
 assign n1407 = ( (~ n314)  &  (~ n350) ) | ( (~ n314)  &  n1473 ) | ( n350  &  n1473 ) ;
 assign n1409 = ( (~ n1565)  &  (~ n2390) ) ;
 assign n1410 = ( (~ n540)  &  n551 ) ;
 assign n1408 = ( n544  &  n1409  &  n1410 ) ;
 assign n1411 = ( (~ n167)  &  n1408 ) | ( (~ n167)  &  (~ n1565)  &  (~ n1566) ) ;
 assign n1415 = ( n540  &  n913  &  (~ n1411) ) | ( n913  &  (~ n1411)  &  (~ n2394) ) ;
 assign n1418 = ( n1897  &  n1473 ) ;
 assign n1417 = ( n1415  &  n1418 ) | ( n1415  &  (~ n2787) ) ;
 assign n1423 = ( n2102  &  n2105 ) | ( (~ n2104)  &  n2105 ) | ( n2102  &  n2107 ) | ( (~ n2104)  &  n2107 ) ;
 assign n1424 = ( n272  &  Ng117 ) | ( (~ n272)  &  (~ Ng117) ) ;
 assign n1422 = ( (~ n1428)  &  (~ n3822) ) | ( n1423  &  n1424  &  (~ n1428) ) ;
 assign n1428 = ( n460 ) | ( (~ Ng2257) ) ;
 assign n1429 = ( n1424 ) | ( n1433 ) | ( n2101 ) | ( n2102 ) | ( (~ n2104) ) | ( n2105 ) | ( n2107 ) | ( n2424 ) ;
 assign n1427 = ( n1428  &  (~ n2429) ) | ( n1429  &  (~ n2429) ) ;
 assign n1432 = ( n2095  &  n2099 ) | ( n2097  &  n2099 ) | ( n2095  &  n2101 ) | ( n2097  &  n2101 ) ;
 assign n1433 = ( (~ n208)  &  n625 ) | ( n208  &  (~ n625) ) ;
 assign n1431 = ( (~ n1428)  &  (~ n3815) ) | ( (~ n1428)  &  n1432  &  n1433 ) ;
 assign n1438 = ( n2108  &  (~ n2119)  &  (~ n2432) ) ;
 assign n1437 = ( n272  &  n1438 ) | ( n1438  &  (~ n1481) ) ;
 assign n1439 = ( n197  &  n1481 ) | ( (~ n197)  &  (~ n1481) ) ;
 assign n1440 = ( (~ n272)  &  (~ n300) ) | ( (~ n272)  &  n1481 ) | ( n300  &  n1481 ) ;
 assign n1442 = ( (~ n1575)  &  (~ n2425) ) ;
 assign n1443 = ( (~ n534)  &  n542 ) ;
 assign n1441 = ( n538  &  n1442  &  n1443 ) ;
 assign n1444 = ( (~ n160)  &  n1441 ) | ( (~ n160)  &  (~ n1575)  &  (~ n1576) ) ;
 assign n1448 = ( n534  &  n908  &  (~ n1444) ) | ( n908  &  (~ n1444)  &  (~ n2429) ) ;
 assign n1451 = ( n1901  &  n1481 ) ;
 assign n1450 = ( n1448  &  n1451 ) | ( n1448  &  (~ n2807) ) ;
 assign n1457 = ( (~ n555) ) | ( n562 ) | ( (~ n567) ) ;
 assign n1455 = ( (~ n414)  &  n1338 ) | ( n1338  &  n1457 ) ;
 assign n1458 = ( n1455  &  n1340 ) ;
 assign n1459 = ( Ng2200  &  (~ n1349) ) ;
 assign n1460 = ( Ng2195  &  (~ n1349) ) ;
 assign n1461 = ( Ng2185  &  (~ n1349) ) ;
 assign n1462 = ( Ng2165  &  (~ n1349) ) ;
 assign n1465 = ( (~ n546) ) | ( n553 ) | ( (~ n560) ) ;
 assign n1463 = ( (~ n364)  &  n1371 ) | ( n1371  &  n1465 ) ;
 assign n1466 = ( n1463  &  n1373 ) ;
 assign n1467 = ( Ng1506  &  (~ n1382) ) ;
 assign n1468 = ( Ng1501  &  (~ n1382) ) ;
 assign n1469 = ( Ng1491  &  (~ n1382) ) ;
 assign n1470 = ( Ng1471  &  (~ n1382) ) ;
 assign n1473 = ( (~ n540) ) | ( n544 ) | ( (~ n551) ) ;
 assign n1471 = ( (~ n314)  &  n1404 ) | ( n1404  &  n1473 ) ;
 assign n1474 = ( n1471  &  n1406 ) ;
 assign n1475 = ( Ng813  &  (~ n1415) ) ;
 assign n1476 = ( Ng809  &  (~ n1415) ) ;
 assign n1477 = ( Ng801  &  (~ n1415) ) ;
 assign n1478 = ( Ng785  &  (~ n1415) ) ;
 assign n1481 = ( (~ n534) ) | ( n538 ) | ( (~ n542) ) ;
 assign n1479 = ( (~ n272)  &  n1437 ) | ( n1437  &  n1481 ) ;
 assign n1482 = ( n1479  &  n1439 ) ;
 assign n1483 = ( Ng125  &  (~ n1448) ) ;
 assign n1484 = ( Ng121  &  (~ n1448) ) ;
 assign n1485 = ( Ng113  &  (~ n1448) ) ;
 assign n1486 = ( Ng97  &  (~ n1448) ) ;
 assign n1488 = ( n497  &  (~ n3824) ) | ( wire1603  &  n497  &  (~ Ng1425) ) ;
 assign n1487 = ( n254  &  n396  &  n431  &  n469  &  n1488  &  (~ n3826) ) ;
 assign n1491 = ( (~ Ng1243)  &  n4034 ) | ( n4032  &  n4034 ) ;
 assign n1490 = ( n1167  &  n1172 ) | ( (~ n1167)  &  (~ n1172) ) ;
 assign n1494 = ( n669 ) | ( (~ n671) ) ;
 assign n1497 = ( (~ n1056) ) | ( n1494 ) ;
 assign n1500 = ( (~ wire1603)  &  (~ Ng1315) ) | ( (~ Ng1315)  &  Ng1422 ) | ( (~ wire1603)  &  Ng1420 ) | ( Ng1422  &  Ng1420 ) ;
 assign n1507 = ( n555  &  n1457 ) | ( n1457  &  (~ n1546) ) | ( n1457  &  (~ n2320) ) ;
 assign n1510 = ( Ng2133  &  Ng2129  &  n1598 ) ;
 assign n1509 = ( n1510  &  Ng2124 ) ;
 assign n1511 = ( n546  &  n1465 ) | ( n1465  &  (~ n1556) ) | ( n1465  &  (~ n2355) ) ;
 assign n1514 = ( Ng1439  &  Ng1435  &  n1605 ) ;
 assign n1513 = ( n1514  &  Ng1430 ) ;
 assign n1515 = ( n540  &  n1473 ) | ( n1473  &  (~ n1566) ) | ( n1473  &  (~ n2390) ) ;
 assign n1518 = ( Ng753  &  Ng749  &  n1612 ) ;
 assign n1517 = ( n1518  &  Ng744 ) ;
 assign n1519 = ( n534  &  n1481 ) | ( n1481  &  (~ n1576) ) | ( n1481  &  (~ n2425) ) ;
 assign n1522 = ( Ng65  &  Ng61  &  n1619 ) ;
 assign n1521 = ( n1522  &  Ng56 ) ;
 assign n1526 = ( n2453 ) | ( n1525 ) ;
 assign n1524 = ( (~ Ng3135) ) | ( n2460 ) ;
 assign n1525 = ( (~ Ng3147) ) | ( n1768 ) ;
 assign n1523 = ( n1526  &  n1524 ) | ( n1526  &  n1525 ) ;
 assign n1529 = ( Ng3120  &  n2497 ) | ( (~ Ng3135)  &  n2497 ) | ( n2497  &  (~ n2954) ) ;
 assign n1527 = ( Ng3147 ) | ( n1768 ) | ( n1524 ) ;
 assign n1530 = ( wire1605  &  (~ Ng8284) ) ;
 assign n1533 = ( n462  &  (~ n3836) ) | ( wire1603  &  n462  &  (~ Ng739) ) ;
 assign n1532 = ( n226  &  n346  &  n381  &  n424  &  n1533  &  (~ n3838) ) ;
 assign n1536 = ( (~ Ng557)  &  n4057 ) | ( n4055  &  n4057 ) ;
 assign n1535 = ( n1153  &  n1158 ) | ( (~ n1153)  &  (~ n1158) ) ;
 assign n1541 = ( (~ n629) ) | ( (~ n1215) ) | ( (~ Ng2257) ) | ( (~ n2324) ) ;
 assign n1538 = ( n629  &  n657 ) | ( n629  &  (~ n1215) ) ;
 assign n1539 = ( (~ n629)  &  n657 ) | ( (~ n629)  &  n1215 ) ;
 assign n1540 = ( n620 ) | ( (~ Ng2257) ) ;
 assign n1537 = ( n1541  &  n1538 ) | ( n1541  &  n1539 ) | ( n1541  &  n1540 ) ;
 assign n1545 = ( n1994 ) | ( n1995 ) | ( n1329 ) | ( n2295 ) | ( n2296 ) | ( n2297 ) ;
 assign n1546 = ( n555 ) | ( (~ n562) ) | ( n567 ) ;
 assign n1542 = ( (~ n1343)  &  n1545 ) | ( (~ n1344)  &  n1545 ) | ( (~ n1343)  &  n1546 ) | ( (~ n1344)  &  n1546 ) ;
 assign n1551 = ( (~ n615) ) | ( (~ n1212) ) | ( (~ Ng2257) ) | ( (~ n2359) ) ;
 assign n1548 = ( n615  &  n652 ) | ( n615  &  (~ n1212) ) ;
 assign n1549 = ( (~ n615)  &  n652 ) | ( (~ n615)  &  n1212 ) ;
 assign n1550 = ( n606 ) | ( (~ Ng2257) ) ;
 assign n1547 = ( n1551  &  n1548 ) | ( n1551  &  n1549 ) | ( n1551  &  n1550 ) ;
 assign n1555 = ( n2027 ) | ( n2028 ) | ( n1362 ) | ( n2330 ) | ( n2331 ) | ( n2332 ) ;
 assign n1556 = ( n546 ) | ( (~ n553) ) | ( n560 ) ;
 assign n1552 = ( (~ n1376)  &  n1555 ) | ( (~ n1377)  &  n1555 ) | ( (~ n1376)  &  n1556 ) | ( (~ n1377)  &  n1556 ) ;
 assign n1561 = ( (~ n601) ) | ( (~ n1209) ) | ( (~ Ng2257) ) | ( (~ n2394) ) ;
 assign n1558 = ( n601  &  n647 ) | ( n601  &  (~ n1209) ) ;
 assign n1559 = ( (~ n601)  &  n647 ) | ( (~ n601)  &  n1209 ) ;
 assign n1560 = ( n592 ) | ( (~ Ng2257) ) ;
 assign n1557 = ( n1561  &  n1558 ) | ( n1561  &  n1559 ) | ( n1561  &  n1560 ) ;
 assign n1565 = ( n2060 ) | ( n2061 ) | ( n1395 ) | ( n2365 ) | ( n2366 ) | ( n2367 ) ;
 assign n1566 = ( n540 ) | ( (~ n544) ) | ( n551 ) ;
 assign n1562 = ( (~ n1409)  &  n1565 ) | ( (~ n1410)  &  n1565 ) | ( (~ n1409)  &  n1566 ) | ( (~ n1410)  &  n1566 ) ;
 assign n1571 = ( (~ n587) ) | ( (~ n1206) ) | ( (~ Ng2257) ) | ( (~ n2429) ) ;
 assign n1568 = ( n587  &  n645 ) | ( n587  &  (~ n1206) ) ;
 assign n1569 = ( (~ n587)  &  n645 ) | ( (~ n587)  &  n1206 ) ;
 assign n1570 = ( n578 ) | ( (~ Ng2257) ) ;
 assign n1567 = ( n1571  &  n1568 ) | ( n1571  &  n1569 ) | ( n1571  &  n1570 ) ;
 assign n1575 = ( n2093 ) | ( n2094 ) | ( n1428 ) | ( n2400 ) | ( n2401 ) | ( n2402 ) ;
 assign n1576 = ( n534 ) | ( (~ n538) ) | ( n542 ) ;
 assign n1572 = ( (~ n1442)  &  n1575 ) | ( (~ n1443)  &  n1575 ) | ( (~ n1442)  &  n1576 ) | ( (~ n1443)  &  n1576 ) ;
 assign n1579 = ( n665 ) | ( (~ n667) ) ;
 assign n1582 = ( (~ n1015) ) | ( n1579 ) ;
 assign n1585 = ( (~ wire1603)  &  (~ Ng1315) ) | ( (~ Ng1315)  &  Ng736 ) | ( (~ wire1603)  &  Ng734 ) | ( Ng736  &  Ng734 ) ;
 assign n1595 = ( n629 ) | ( (~ n657) ) | ( n1215 ) ;
 assign n1593 = ( (~ n657)  &  (~ n1540)  &  n1595 ) | ( n1216  &  (~ n1540)  &  n1595 ) ;
 assign n1598 = ( Ng2142  &  Ng2138  &  n1796 ) ;
 assign n1597 = ( n1598  &  Ng2133 ) ;
 assign n1602 = ( n615 ) | ( (~ n652) ) | ( n1212 ) ;
 assign n1600 = ( (~ n652)  &  (~ n1550)  &  n1602 ) | ( n1213  &  (~ n1550)  &  n1602 ) ;
 assign n1605 = ( Ng1448  &  Ng1444  &  n1806 ) ;
 assign n1604 = ( n1605  &  Ng1439 ) ;
 assign n1609 = ( n601 ) | ( (~ n647) ) | ( n1209 ) ;
 assign n1607 = ( (~ n647)  &  (~ n1560)  &  n1609 ) | ( n1210  &  (~ n1560)  &  n1609 ) ;
 assign n1612 = ( Ng762  &  Ng758  &  n1816 ) ;
 assign n1611 = ( n1612  &  Ng753 ) ;
 assign n1616 = ( n587 ) | ( (~ n645) ) | ( n1206 ) ;
 assign n1614 = ( (~ n645)  &  (~ n1570)  &  n1616 ) | ( n1207  &  (~ n1570)  &  n1616 ) ;
 assign n1619 = ( Ng74  &  Ng70  &  n1826 ) ;
 assign n1618 = ( n1619  &  Ng65 ) ;
 assign n1620 = ( (~ wire1521)  &  n1523 ) ;
 assign n1621 = ( n1527  &  (~ Ng3105) ) | ( n1527  &  n2521 ) | ( (~ Ng3105)  &  Ng3128 ) | ( n2521  &  Ng3128 ) ;
 assign n1622 = ( (~ Ng3104)  &  (~ Ng3103) ) | ( (~ Ng3104)  &  n2519 ) | ( (~ Ng3103)  &  n2520 ) | ( n2519  &  n2520 ) ;
 assign n1623 = ( n2515  &  n2517 ) | ( (~ Ng3101)  &  n2517 ) | ( n2515  &  (~ Ng3102) ) | ( (~ Ng3101)  &  (~ Ng3102) ) ;
 assign n1624 = ( n2510  &  n2512 ) | ( (~ Ng3099)  &  n2512 ) | ( n2510  &  (~ Ng3100) ) | ( (~ Ng3099)  &  (~ Ng3100) ) ;
 assign n1625 = ( n2506  &  n2508 ) | ( (~ Ng3097)  &  n2508 ) | ( n2506  &  (~ Ng3098) ) | ( (~ Ng3097)  &  (~ Ng3098) ) ;
 assign n1626 = ( (~ Ng3108)  &  (~ Ng3107) ) | ( (~ Ng3108)  &  n2502 ) | ( (~ Ng3107)  &  n2504 ) | ( n2502  &  n2504 ) ;
 assign n1627 = ( (~ Ng3106)  &  n2497 ) | ( n2497  &  n2501 ) | ( (~ Ng3106)  &  (~ n4878) ) | ( n2501  &  (~ n4878) ) ;
 assign n1629 = ( Ng2753  &  n2523 ) ;
 assign n1628 = ( Ng2760  &  n1629 ) ;
 assign n1630 = ( n103  &  (~ n112) ) | ( (~ n112)  &  (~ n599) ) | ( n103  &  (~ n623) ) | ( (~ n599)  &  (~ n623) ) ;
 assign n1634 = ( n599  &  (~ n3850) ) | ( n109  &  n599  &  (~ n623) ) ;
 assign n1636 = ( n112  &  (~ n3848) ) | ( n103  &  n112  &  (~ n611) ) ;
 assign n1640 = ( n623  &  n611 ) ;
 assign n1639 = ( (~ n599)  &  n1636 ) | ( n94  &  (~ n599)  &  n1640 ) ;
 assign n1641 = ( (~ n112)  &  n1634 ) | ( (~ n112)  &  (~ n632)  &  (~ n1654) ) ;
 assign n1646 = ( n94 ) | ( n109 ) | ( (~ n623) ) ;
 assign n1644 = ( (~ n103)  &  n1646 ) | ( n109  &  (~ n623)  &  n1646 ) ;
 assign n1647 = ( n112  &  n623 ) | ( n623  &  (~ n632) ) ;
 assign n1648 = ( n103  &  (~ n632) ) | ( n103  &  (~ n109)  &  n1640 ) ;
 assign n1650 = ( n94  &  (~ n1648) ) | ( n599  &  (~ n1648) ) | ( n632  &  (~ n1648) ) ;
 assign n1653 = ( n112  &  (~ n611) ) | ( (~ n112)  &  n623 ) | ( (~ n611)  &  n623 ) ;
 assign n1654 = ( n103 ) | ( n109 ) ;
 assign n1652 = ( (~ n94)  &  n1653 ) | ( n1647  &  n1653 ) | ( (~ n94)  &  n1654 ) | ( n1647  &  n1654 ) ;
 assign n1657 = ( n611 ) | ( n1644 ) | ( n112 ) ;
 assign n1658 = ( n599  &  n1652 ) | ( (~ n599)  &  (~ n3000) ) | ( n1652  &  (~ n3000) ) ;
 assign n1656 = ( (~ n112)  &  n1657  &  n1658 ) | ( n1650  &  n1657  &  n1658 ) ;
 assign n1661 = ( Ng16474 ) | ( (~ Ng185) ) | ( (~ Ng2616) ) ;
 assign n1662 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1605)  &  (~ Ng2673) ) | ( (~ wire1603)  &  (~ Ng2670) ) | ( (~ Ng2673)  &  (~ Ng2670) ) ;
 assign n1659 = ( (~ Ng1315)  &  n1661  &  n1662 ) | ( n1661  &  n1662  &  (~ Ng2676) ) ;
 assign n1664 = ( Ng2059  &  n2551 ) ;
 assign n1663 = ( Ng2066  &  n1664 ) ;
 assign n1665 = ( n91  &  (~ n106) ) | ( (~ n106)  &  (~ n585) ) | ( n91  &  (~ n609) ) | ( (~ n585)  &  (~ n609) ) ;
 assign n1669 = ( n585  &  (~ n3853) ) | ( n100  &  n585  &  (~ n609) ) ;
 assign n1671 = ( n106  &  (~ n3851) ) | ( n91  &  n106  &  (~ n597) ) ;
 assign n1675 = ( n609  &  n597 ) ;
 assign n1674 = ( (~ n585)  &  n1671 ) | ( n82  &  (~ n585)  &  n1675 ) ;
 assign n1676 = ( (~ n106)  &  n1669 ) | ( (~ n106)  &  (~ n618)  &  (~ n1689) ) ;
 assign n1681 = ( n82 ) | ( n100 ) | ( (~ n609) ) ;
 assign n1679 = ( (~ n91)  &  n1681 ) | ( n100  &  (~ n609)  &  n1681 ) ;
 assign n1682 = ( n106  &  n609 ) | ( n609  &  (~ n618) ) ;
 assign n1683 = ( n91  &  (~ n618) ) | ( n91  &  (~ n100)  &  n1675 ) ;
 assign n1685 = ( n82  &  (~ n1683) ) | ( n585  &  (~ n1683) ) | ( n618  &  (~ n1683) ) ;
 assign n1688 = ( n106  &  (~ n597) ) | ( (~ n106)  &  n609 ) | ( (~ n597)  &  n609 ) ;
 assign n1689 = ( n91 ) | ( n100 ) ;
 assign n1687 = ( (~ n82)  &  n1688 ) | ( n1682  &  n1688 ) | ( (~ n82)  &  n1689 ) | ( n1682  &  n1689 ) ;
 assign n1692 = ( n597 ) | ( n1679 ) | ( n106 ) ;
 assign n1693 = ( n585  &  n1687 ) | ( (~ n585)  &  (~ n3013) ) | ( n1687  &  (~ n3013) ) ;
 assign n1691 = ( (~ n106)  &  n1692  &  n1693 ) | ( n1685  &  n1692  &  n1693 ) ;
 assign n1696 = ( Ng16472 ) | ( (~ Ng185) ) | ( (~ Ng1922) ) ;
 assign n1697 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1605)  &  (~ Ng1979) ) | ( (~ wire1603)  &  (~ Ng1976) ) | ( (~ Ng1979)  &  (~ Ng1976) ) ;
 assign n1694 = ( (~ Ng1315)  &  n1696  &  n1697 ) | ( n1696  &  n1697  &  (~ Ng1982) ) ;
 assign n1699 = ( Ng1365  &  n2575 ) ;
 assign n1698 = ( Ng1372  &  n1699 ) ;
 assign n1700 = ( n79  &  (~ n97) ) | ( (~ n97)  &  (~ n576) ) | ( n79  &  (~ n595) ) | ( (~ n576)  &  (~ n595) ) ;
 assign n1704 = ( n576  &  (~ n3856) ) | ( n88  &  n576  &  (~ n595) ) ;
 assign n1706 = ( n97  &  (~ n3854) ) | ( n79  &  n97  &  (~ n583) ) ;
 assign n1710 = ( n595  &  n583 ) ;
 assign n1709 = ( (~ n576)  &  n1706 ) | ( n73  &  (~ n576)  &  n1710 ) ;
 assign n1711 = ( (~ n97)  &  n1704 ) | ( (~ n97)  &  (~ n604)  &  (~ n1724) ) ;
 assign n1716 = ( n73 ) | ( n88 ) | ( (~ n595) ) ;
 assign n1714 = ( (~ n79)  &  n1716 ) | ( n88  &  (~ n595)  &  n1716 ) ;
 assign n1717 = ( n97  &  n595 ) | ( n595  &  (~ n604) ) ;
 assign n1718 = ( n79  &  (~ n604) ) | ( n79  &  (~ n88)  &  n1710 ) ;
 assign n1720 = ( n73  &  (~ n1718) ) | ( n576  &  (~ n1718) ) | ( n604  &  (~ n1718) ) ;
 assign n1723 = ( n97  &  (~ n583) ) | ( (~ n97)  &  n595 ) | ( (~ n583)  &  n595 ) ;
 assign n1724 = ( n79 ) | ( n88 ) ;
 assign n1722 = ( (~ n73)  &  n1723 ) | ( n1717  &  n1723 ) | ( (~ n73)  &  n1724 ) | ( n1717  &  n1724 ) ;
 assign n1727 = ( n583 ) | ( n1714 ) | ( n97 ) ;
 assign n1728 = ( n576  &  n1722 ) | ( (~ n576)  &  (~ n3026) ) | ( n1722  &  (~ n3026) ) ;
 assign n1726 = ( (~ n97)  &  n1727  &  n1728 ) | ( n1720  &  n1727  &  n1728 ) ;
 assign n1731 = ( Ng16470 ) | ( (~ Ng185) ) | ( (~ Ng1228) ) ;
 assign n1732 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1605)  &  (~ Ng1285) ) | ( (~ wire1603)  &  (~ Ng1282) ) | ( (~ Ng1285)  &  (~ Ng1282) ) ;
 assign n1729 = ( (~ Ng1315)  &  n1731  &  n1732 ) | ( n1731  &  n1732  &  (~ Ng1288) ) ;
 assign n1734 = ( Ng679  &  n2599 ) ;
 assign n1733 = ( Ng686  &  n1734 ) ;
 assign n1735 = ( n70  &  (~ n85) ) | ( (~ n85)  &  (~ n572) ) | ( n70  &  (~ n581) ) | ( (~ n572)  &  (~ n581) ) ;
 assign n1739 = ( n572  &  (~ n3859) ) | ( n76  &  n572  &  (~ n581) ) ;
 assign n1741 = ( n85  &  (~ n3857) ) | ( n70  &  n85  &  (~ n574) ) ;
 assign n1745 = ( n581  &  n574 ) ;
 assign n1744 = ( (~ n572)  &  n1741 ) | ( n66  &  (~ n572)  &  n1745 ) ;
 assign n1746 = ( (~ n85)  &  n1739 ) | ( (~ n85)  &  (~ n590)  &  (~ n1759) ) ;
 assign n1751 = ( n66 ) | ( n76 ) | ( (~ n581) ) ;
 assign n1749 = ( (~ n70)  &  n1751 ) | ( n76  &  (~ n581)  &  n1751 ) ;
 assign n1752 = ( n85  &  n581 ) | ( n581  &  (~ n590) ) ;
 assign n1753 = ( n70  &  (~ n590) ) | ( n70  &  (~ n76)  &  n1745 ) ;
 assign n1755 = ( n66  &  (~ n1753) ) | ( n572  &  (~ n1753) ) | ( n590  &  (~ n1753) ) ;
 assign n1758 = ( n85  &  (~ n574) ) | ( (~ n85)  &  n581 ) | ( (~ n574)  &  n581 ) ;
 assign n1759 = ( n70 ) | ( n76 ) ;
 assign n1757 = ( (~ n66)  &  n1758 ) | ( n1752  &  n1758 ) | ( (~ n66)  &  n1759 ) | ( n1752  &  n1759 ) ;
 assign n1762 = ( n574 ) | ( n1749 ) | ( n85 ) ;
 assign n1763 = ( n572  &  n1757 ) | ( (~ n572)  &  (~ n3039) ) | ( n1757  &  (~ n3039) ) ;
 assign n1761 = ( (~ n85)  &  n1762  &  n1763 ) | ( n1755  &  n1762  &  n1763 ) ;
 assign n1766 = ( Ng16468 ) | ( (~ Ng185) ) | ( (~ Ng542) ) ;
 assign n1767 = ( (~ wire1603)  &  (~ wire1605) ) | ( (~ wire1605)  &  (~ Ng599) ) | ( (~ wire1603)  &  (~ Ng596) ) | ( (~ Ng599)  &  (~ Ng596) ) ;
 assign n1764 = ( (~ Ng1315)  &  n1766  &  n1767 ) | ( n1766  &  n1767  &  (~ Ng602) ) ;
 assign n1768 = ( Ng3126 ) | ( Ng3191 ) | ( Ng3126 ) | ( Ng3110 ) ;
 assign n1769 = ( n1526  &  n1527 ) ;
 assign n1771 = ( n2506  &  n2510 ) | ( n2506  &  (~ Ng3161) ) | ( n2510  &  (~ Ng3155) ) | ( (~ Ng3161)  &  (~ Ng3155) ) ;
 assign n1772 = ( n2508  &  n2512 ) | ( n2508  &  (~ Ng3164) ) | ( n2512  &  (~ Ng3158) ) | ( (~ Ng3164)  &  (~ Ng3158) ) ;
 assign n1773 = ( n2515  &  n2517 ) | ( n2517  &  (~ Ng3167) ) | ( n2515  &  (~ Ng3170) ) | ( (~ Ng3167)  &  (~ Ng3170) ) ;
 assign n1774 = ( n2520  &  n2521 ) | ( n2521  &  (~ Ng3176) ) | ( n2520  &  (~ Ng3179) ) | ( (~ Ng3176)  &  (~ Ng3179) ) ;
 assign n1775 = ( n2519 ) | ( (~ Ng3173) ) ;
 assign n1776 = ( n2501  &  n2502 ) | ( n2501  &  (~ Ng3185) ) | ( n2502  &  (~ Ng3182) ) | ( (~ Ng3185)  &  (~ Ng3182) ) ;
 assign n1777 = ( n1769  &  n2504 ) | ( (~ Ng3135)  &  n2504 ) | ( n1769  &  (~ Ng3088) ) | ( (~ Ng3135)  &  (~ Ng3088) ) ;
 assign n1770 = ( (~ wire1521)  &  n1771  &  n1772  &  n1773  &  n1774  &  n1775  &  n1776  &  n1777 ) ;
 assign n1779 = ( n2502  &  n2504 ) | ( n2504  &  (~ Ng3095) ) | ( n2502  &  (~ Ng3096) ) | ( (~ Ng3095)  &  (~ Ng3096) ) ;
 assign n1780 = ( n2501  &  n2521 ) | ( n2501  &  (~ Ng3093) ) | ( n2521  &  (~ Ng3094) ) | ( (~ Ng3093)  &  (~ Ng3094) ) ;
 assign n1781 = ( n2519  &  n2520 ) | ( n2520  &  (~ Ng3091) ) | ( n2519  &  (~ Ng3092) ) | ( (~ Ng3091)  &  (~ Ng3092) ) ;
 assign n1782 = ( n2515  &  n2517 ) | ( n2517  &  (~ Ng3086) ) | ( n2515  &  (~ Ng3087) ) | ( (~ Ng3086)  &  (~ Ng3087) ) ;
 assign n1783 = ( n2510  &  n2512 ) | ( n2512  &  (~ Ng3084) ) | ( n2510  &  (~ Ng3085) ) | ( (~ Ng3084)  &  (~ Ng3085) ) ;
 assign n1784 = ( n2506  &  n2508 ) | ( n2508  &  (~ Ng3210) ) | ( n2506  &  (~ Ng3211) ) | ( (~ Ng3210)  &  (~ Ng3211) ) ;
 assign n1785 = ( (~ Ng3120)  &  n3860 ) | ( n1523  &  n1527  &  n3860 ) ;
 assign n1778 = ( (~ wire1521)  &  n1779  &  n1780  &  n1781  &  n1782  &  n1783  &  n1784  &  n1785 ) ;
 assign n1789 = ( Ng2195  &  Ng2200  &  Ng2185  &  Ng2190  &  Ng2175  &  Ng2180  &  Ng2165  &  Ng2170 ) ;
 assign n1786 = ( n1789  &  (~ n3861) ) | ( wire1594  &  n1789  &  (~ Ng2255) ) ;
 assign n1791 = ( n455  &  (~ n488) ) | ( n455  &  (~ n1786) ) ;
 assign n1792 = ( (~ n455)  &  n488 ) | ( (~ n455)  &  n1786 ) ;
 assign n1790 = ( (~ Ng2257) ) | ( n1791 ) | ( n1792 ) ;
 assign n1796 = ( Ng2151  &  Ng2147  &  n1873 ) ;
 assign n1795 = ( n1796  &  Ng2142 ) ;
 assign n1800 = ( Ng1501  &  Ng1506  &  Ng1491  &  Ng1496  &  Ng1481  &  Ng1486  &  Ng1471  &  Ng1476 ) ;
 assign n1797 = ( n1800  &  (~ n3862) ) | ( wire1594  &  n1800  &  (~ Ng1561) ) ;
 assign n1802 = ( n405  &  (~ n443) ) | ( n405  &  (~ n1797) ) ;
 assign n1803 = ( (~ n405)  &  n443 ) | ( (~ n405)  &  n1797 ) ;
 assign n1801 = ( (~ Ng2257) ) | ( n1802 ) | ( n1803 ) ;
 assign n1806 = ( Ng1457  &  Ng1453  &  n1877 ) ;
 assign n1805 = ( n1806  &  Ng1448 ) ;
 assign n1810 = ( Ng809  &  Ng813  &  Ng801  &  Ng805  &  Ng793  &  Ng797  &  Ng785  &  Ng789 ) ;
 assign n1807 = ( n1810  &  (~ n3863) ) | ( wire1594  &  n1810  &  (~ Ng867) ) ;
 assign n1812 = ( n355  &  (~ n393) ) | ( n355  &  (~ n1807) ) ;
 assign n1813 = ( (~ n355)  &  n393 ) | ( (~ n355)  &  n1807 ) ;
 assign n1811 = ( (~ Ng2257) ) | ( n1812 ) | ( n1813 ) ;
 assign n1816 = ( Ng771  &  Ng767  &  n1881 ) ;
 assign n1815 = ( n1816  &  Ng762 ) ;
 assign n1820 = ( Ng121  &  Ng125  &  Ng113  &  Ng117  &  Ng105  &  Ng109  &  Ng97  &  Ng101 ) ;
 assign n1817 = ( n1820  &  (~ n3864) ) | ( wire1594  &  n1820  &  (~ Ng179) ) ;
 assign n1822 = ( n305  &  (~ n343) ) | ( n305  &  (~ n1817) ) ;
 assign n1823 = ( (~ n305)  &  n343 ) | ( (~ n305)  &  n1817 ) ;
 assign n1821 = ( (~ Ng2257) ) | ( n1822 ) | ( n1823 ) ;
 assign n1826 = ( Ng83  &  Ng79  &  n1885 ) ;
 assign n1825 = ( n1826  &  Ng74 ) ;
 assign n1830 = ( (~ n124) ) | ( n569 ) | ( (~ Ng2584) ) ;
 assign n1834 = ( Pg3229 ) | ( n611 ) | ( (~ n623) ) ;
 assign n1831 = ( (~ Pg3229)  &  n1834  &  (~ n4158) ) | ( n632  &  n1834  &  (~ n4158) ) ;
 assign n1837 = ( Pg3229 ) | ( n486 ) | ( (~ n509) ) ;
 assign n1835 = ( (~ Pg3229)  &  n1837  &  (~ n4181) ) | ( n524  &  n1837  &  (~ n4181) ) ;
 assign n1840 = ( (~ n121) ) | ( n564 ) | ( (~ Ng1890) ) ;
 assign n1843 = ( Pg3229 ) | ( n597 ) | ( (~ n609) ) ;
 assign n1841 = ( (~ Pg3229)  &  n1843  &  (~ n4205) ) | ( n618  &  n1843  &  (~ n4205) ) ;
 assign n1846 = ( Pg3229 ) | ( n441 ) | ( (~ n474) ) ;
 assign n1844 = ( (~ Pg3229)  &  n1846  &  (~ n4228) ) | ( n502  &  n1846  &  (~ n4228) ) ;
 assign n1849 = ( (~ n118) ) | ( n557 ) | ( (~ Ng1196) ) ;
 assign n1852 = ( Pg3229 ) | ( n583 ) | ( (~ n595) ) ;
 assign n1850 = ( (~ Pg3229)  &  n1852  &  (~ n4252) ) | ( n604  &  n1852  &  (~ n4252) ) ;
 assign n1855 = ( Pg3229 ) | ( n391 ) | ( (~ n429) ) ;
 assign n1853 = ( (~ Pg3229)  &  n1855  &  (~ n4275) ) | ( n467  &  n1855  &  (~ n4275) ) ;
 assign n1858 = ( (~ n115) ) | ( n548 ) | ( (~ Ng510) ) ;
 assign n1861 = ( Pg3229 ) | ( n574 ) | ( (~ n581) ) ;
 assign n1859 = ( (~ Pg3229)  &  n1861  &  (~ n4299) ) | ( n590  &  n1861  &  (~ n4299) ) ;
 assign n1864 = ( Pg3229 ) | ( n341 ) | ( (~ n379) ) ;
 assign n1862 = ( (~ Pg3229)  &  n1864  &  (~ n4322) ) | ( n422  &  n1864  &  (~ n4322) ) ;
 assign n1867 = ( (~ Ng3013) ) | ( n2695 ) ;
 assign n1865 = ( n1867 ) | ( (~ Ng3010) ) ;
 assign n1869 = ( Ng2903  &  n2699 ) ;
 assign n1868 = ( Ng2900  &  n1869 ) ;
 assign n1871 = ( Ng2734  &  Ng2720  &  n1914 ) ;
 assign n1870 = ( n1871  &  Ng2746 ) ;
 assign n1873 = ( (~ n1916)  &  Ng2160  &  Ng2156 ) ;
 assign n1872 = ( n1873  &  Ng2151 ) ;
 assign n1875 = ( Ng2040  &  Ng2026  &  n1919 ) ;
 assign n1874 = ( n1875  &  Ng2052 ) ;
 assign n1877 = ( (~ n1916)  &  Ng1466  &  Ng1462 ) ;
 assign n1876 = ( n1877  &  Ng1457 ) ;
 assign n1879 = ( Ng1346  &  Ng1332  &  n1923 ) ;
 assign n1878 = ( n1879  &  Ng1358 ) ;
 assign n1881 = ( (~ n1916)  &  Ng780  &  Ng776 ) ;
 assign n1880 = ( n1881  &  Ng771 ) ;
 assign n1883 = ( Ng660  &  Ng646  &  n1927 ) ;
 assign n1882 = ( n1883  &  Ng672 ) ;
 assign n1885 = ( (~ n1916)  &  Ng92  &  Ng88 ) ;
 assign n1884 = ( n1885  &  Ng83 ) ;
 assign n1886 = ( (~ n721) ) | ( (~ n733) ) | ( n2145 ) | ( n2146 ) | ( n2147 ) | ( n2148 ) ;
 assign n1887 = ( n2152 ) | ( n2153 ) | ( n2154 ) | ( n2149 ) | ( n2150 ) | ( n2151 ) ;
 assign n1889 = ( (~ n555) ) | ( (~ n562) ) | ( (~ n567) ) ;
 assign Ng27229 = ( n1886  &  n1889 ) | ( n1887  &  n1889 ) | ( n1886  &  (~ n2326) ) | ( n1887  &  (~ n2326) ) ;
 assign n1890 = ( (~ n721) ) | ( (~ n730) ) | ( n2156 ) | ( n2157 ) | ( n2158 ) | ( n2159 ) ;
 assign n1891 = ( n2163 ) | ( n2164 ) | ( n2165 ) | ( n2160 ) | ( n2161 ) | ( n2162 ) ;
 assign n1893 = ( (~ n546) ) | ( (~ n553) ) | ( (~ n560) ) ;
 assign Ng27220 = ( n1890  &  n1893 ) | ( n1891  &  n1893 ) | ( n1890  &  (~ n2361) ) | ( n1891  &  (~ n2361) ) ;
 assign n1894 = ( (~ n721) ) | ( (~ n726) ) | ( n2167 ) | ( n2168 ) | ( n2169 ) | ( n2170 ) ;
 assign n1895 = ( n2174 ) | ( n2175 ) | ( n2176 ) | ( n2171 ) | ( n2172 ) | ( n2173 ) ;
 assign n1897 = ( (~ n540) ) | ( (~ n544) ) | ( (~ n551) ) ;
 assign Ng27199 = ( n1894  &  n1897 ) | ( n1895  &  n1897 ) | ( n1894  &  (~ n2396) ) | ( n1895  &  (~ n2396) ) ;
 assign n1898 = ( (~ n722) ) | ( (~ n721) ) | ( n2178 ) | ( n2179 ) | ( n2180 ) | ( n2181 ) ;
 assign n1899 = ( n2185 ) | ( n2186 ) | ( n2187 ) | ( n2182 ) | ( n2183 ) | ( n2184 ) ;
 assign n1901 = ( (~ n534) ) | ( (~ n538) ) | ( (~ n542) ) ;
 assign Ng27190 = ( n1898  &  n1901 ) | ( n1899  &  n1901 ) | ( n1898  &  (~ n2431) ) | ( n1899  &  (~ n2431) ) ;
 assign n1902 = ( Ng3032  &  Ng3018  &  (~ Ng3036)  &  (~ Ng3028) ) ;
 assign n1905 = ( n1936 ) | ( Pg3234 ) ;
 assign n1907 = ( Ng3028  &  Ng3018  &  n1936 ) ;
 assign n1906 = ( n1907  &  Ng3036 ) ;
 assign n1908 = ( Ng2912  &  Ng2920  &  (~ Ng2924)  &  (~ Ng2917) ) ;
 assign n1912 = ( Ng2912  &  Ng2917  &  n1938 ) ;
 assign n1911 = ( n1912  &  Ng2924 ) ;
 assign n1914 = ( Ng2727  &  Ng2707  &  n1940 ) ;
 assign n1913 = ( n1914  &  Ng2720 ) ;
 assign n1916 = ( (~ Ng853) ) | ( (~ n721) ) ;
 assign n1915 = ( n1916 ) | ( (~ Ng2160) ) ;
 assign n1919 = ( Ng2033  &  Ng2013  &  n1942 ) ;
 assign n1918 = ( n1919  &  Ng2026 ) ;
 assign n1920 = ( n1916 ) | ( (~ Ng1466) ) ;
 assign n1923 = ( Ng1339  &  Ng1319  &  n1944 ) ;
 assign n1922 = ( n1923  &  Ng1332 ) ;
 assign n1924 = ( n1916 ) | ( (~ Ng780) ) ;
 assign n1927 = ( Ng653  &  Ng633  &  n1946 ) ;
 assign n1926 = ( n1927  &  Ng646 ) ;
 assign n1928 = ( n1916 ) | ( (~ Ng92) ) ;
 assign n1930 = ( (~ n2694) ) | ( (~ Ng3006) ) ;
 assign n1934 = ( Ng13457  &  Ng2888  &  Ng2883 ) ;
 assign n1933 = ( n1934  &  Ng2896 ) ;
 assign n1936 = ( n2524  &  Ng13475 ) ;
 assign n1935 = ( n1936  &  Ng3018 ) ;
 assign n1938 = ( Ng13457  &  (~ Ng2900)  &  (~ Ng2896)  &  (~ Ng2883)  &  Ng2892  &  Ng2903  &  Ng2908  &  Ng2888 ) ;
 assign n1937 = ( n1938  &  Ng2912 ) ;
 assign n1940 = ( Ng1315  &  (~ Ng2733)  &  Ng2714 ) ;
 assign n1939 = ( n1940  &  Ng2707 ) ;
 assign n1942 = ( Ng1315  &  (~ Ng2039)  &  Ng2020 ) ;
 assign n1941 = ( n1942  &  Ng2013 ) ;
 assign n1944 = ( Ng1315  &  (~ Ng1345)  &  Ng1326 ) ;
 assign n1943 = ( n1944  &  Ng1319 ) ;
 assign n1946 = ( Ng1315  &  (~ Ng659)  &  Ng640 ) ;
 assign n1945 = ( n1946  &  Ng633 ) ;
 assign n1947 = ( Ng2883  &  Ng13457 ) ;
 assign n1948 = ( (~ Ng1315) ) | ( Ng2733 ) ;
 assign n1951 = ( (~ Ng1315) ) | ( n1949 ) ;
 assign n1949 = ( Ng1315  &  n2547 ) ;
 assign n1952 = ( (~ Ng1315) ) | ( Ng2039 ) ;
 assign n1954 = ( (~ Ng1315) ) | ( Ng1345 ) ;
 assign n1956 = ( (~ Ng1315) ) | ( Ng659 ) ;
 assign n1960 = ( (~ Ng1315) ) | ( n1958 ) ;
 assign n1958 = ( n4869  &  Ng1315 ) ;
 assign n1966 = ( n177  &  (~ n1323)  &  n1328 ) | ( (~ n1323)  &  n1328  &  (~ n1343) ) ;
 assign n1968 = ( n173  &  (~ n1356)  &  n1361 ) | ( (~ n1356)  &  n1361  &  (~ n1376) ) ;
 assign n1970 = ( n167  &  (~ n1389)  &  n1394 ) | ( (~ n1389)  &  n1394  &  (~ n1409) ) ;
 assign n1972 = ( n160  &  (~ n1422)  &  n1427 ) | ( (~ n1422)  &  n1427  &  (~ n1442) ) ;
 assign n1976 = ( (~ Ng185) ) | ( (~ Ng3139) ) ;
 assign n1974 = ( n1976  &  Ng3139  &  (~ n2455) ) | ( n1976  &  (~ n2455)  &  (~ n4878) ) ;
 assign n1978 = ( (~ Pg3234)  &  n1905 ) | ( (~ Pg3234)  &  (~ n2142) ) ;
 assign Ng27238 = ( (~ n1978) ) ;
 assign n1988 = ( n293  &  Ng2195 ) | ( (~ n293)  &  (~ Ng2195) ) ;
 assign n1989 = ( n448  &  Ng2170 ) | ( (~ n448)  &  (~ Ng2170) ) ;
 assign n1990 = ( n219  &  Ng2180 ) | ( (~ n219)  &  (~ Ng2180) ) ;
 assign n1991 = ( n204  &  Ng2175 ) | ( (~ n204)  &  (~ Ng2175) ) ;
 assign n1992 = ( n326  &  Ng2200 ) | ( (~ n326)  &  (~ Ng2200) ) ;
 assign n1993 = ( n263  &  Ng2190 ) | ( (~ n263)  &  (~ Ng2190) ) ;
 assign n1994 = ( n240  &  Ng2185 ) | ( (~ n240)  &  (~ Ng2185) ) ;
 assign n1995 = ( n410  &  Ng2165 ) | ( (~ n410)  &  (~ Ng2165) ) ;
 assign n1996 = ( n506  &  Ng2175 ) | ( (~ n506)  &  (~ Ng2175) ) ;
 assign n1998 = ( n480  &  Ng2165 ) | ( (~ n480)  &  (~ Ng2165) ) ;
 assign n2000 = ( n265  &  Ng2195 ) | ( (~ n265)  &  (~ Ng2195) ) ;
 assign n2002 = ( n521  &  Ng2185 ) | ( (~ n521)  &  (~ Ng2185) ) ;
 assign n2003 = ( n371  &  Ng2180 ) | ( (~ n371)  &  (~ Ng2180) ) ;
 assign n2005 = ( n483  &  n640 ) | ( (~ n483)  &  (~ n640) ) ;
 assign n2006 = ( n450  &  Ng2200 ) | ( (~ n450)  &  (~ Ng2200) ) ;
 assign n2008 = ( n328  &  Ng2170 ) | ( (~ n328)  &  (~ Ng2170) ) ;
 assign n2009 = ( n521  &  n1457 ) | ( (~ n521)  &  (~ n1457) ) ;
 assign n2011 = ( (~ n480)  &  n1457 ) | ( n480  &  (~ n1457) ) ;
 assign n2012 = ( (~ n328)  &  n1457 ) | ( n328  &  (~ n1457) ) ;
 assign n2014 = ( (~ n506)  &  n1457 ) | ( n506  &  (~ n1457) ) ;
 assign n2015 = ( (~ n371)  &  n1457 ) | ( n371  &  (~ n1457) ) ;
 assign n2017 = ( n2014 ) | ( n2020 ) ;
 assign n2018 = ( n1352 ) | ( n2011 ) ;
 assign n2020 = ( n2012 ) | ( n2018 ) ;
 assign n2021 = ( n193  &  Ng1481 ) | ( (~ n193)  &  (~ Ng1481) ) ;
 assign n2022 = ( n202  &  Ng1486 ) | ( (~ n202)  &  (~ Ng1486) ) ;
 assign n2023 = ( n360  &  Ng1471 ) | ( (~ n360)  &  (~ Ng1471) ) ;
 assign n2024 = ( n217  &  Ng1491 ) | ( (~ n217)  &  (~ Ng1491) ) ;
 assign n2025 = ( n398  &  Ng1476 ) | ( (~ n398)  &  (~ Ng1476) ) ;
 assign n2026 = ( n235  &  Ng1496 ) | ( (~ n235)  &  (~ Ng1496) ) ;
 assign n2027 = ( n284  &  Ng1506 ) | ( (~ n284)  &  (~ Ng1506) ) ;
 assign n2028 = ( n258  &  Ng1501 ) | ( (~ n258)  &  (~ Ng1501) ) ;
 assign n2029 = ( n471  &  Ng1481 ) | ( (~ n471)  &  (~ Ng1481) ) ;
 assign n2031 = ( n435  &  Ng1471 ) | ( (~ n435)  &  (~ Ng1471) ) ;
 assign n2033 = ( n237  &  Ng1501 ) | ( (~ n237)  &  (~ Ng1501) ) ;
 assign n2035 = ( n499  &  Ng1491 ) | ( (~ n499)  &  (~ Ng1491) ) ;
 assign n2036 = ( n321  &  Ng1486 ) | ( (~ n321)  &  (~ Ng1486) ) ;
 assign n2038 = ( n438  &  n636 ) | ( (~ n438)  &  (~ n636) ) ;
 assign n2039 = ( n400  &  Ng1506 ) | ( (~ n400)  &  (~ Ng1506) ) ;
 assign n2041 = ( n286  &  Ng1476 ) | ( (~ n286)  &  (~ Ng1476) ) ;
 assign n2042 = ( n499  &  n1465 ) | ( (~ n499)  &  (~ n1465) ) ;
 assign n2044 = ( (~ n435)  &  n1465 ) | ( n435  &  (~ n1465) ) ;
 assign n2045 = ( (~ n286)  &  n1465 ) | ( n286  &  (~ n1465) ) ;
 assign n2047 = ( (~ n471)  &  n1465 ) | ( n471  &  (~ n1465) ) ;
 assign n2048 = ( (~ n321)  &  n1465 ) | ( n321  &  (~ n1465) ) ;
 assign n2050 = ( n2047 ) | ( n2053 ) ;
 assign n2051 = ( n1385 ) | ( n2044 ) ;
 assign n2053 = ( n2045 ) | ( n2051 ) ;
 assign n2054 = ( n186  &  Ng793 ) | ( (~ n186)  &  (~ Ng793) ) ;
 assign n2055 = ( n348  &  Ng789 ) | ( (~ n348)  &  (~ Ng789) ) ;
 assign n2056 = ( n249  &  Ng813 ) | ( (~ n249)  &  (~ Ng813) ) ;
 assign n2057 = ( n191  &  Ng797 ) | ( (~ n191)  &  (~ Ng797) ) ;
 assign n2058 = ( n230  &  Ng809 ) | ( (~ n230)  &  (~ Ng809) ) ;
 assign n2059 = ( n212  &  Ng805 ) | ( (~ n212)  &  (~ Ng805) ) ;
 assign n2060 = ( n200  &  Ng801 ) | ( (~ n200)  &  (~ Ng801) ) ;
 assign n2061 = ( n310  &  Ng785 ) | ( (~ n310)  &  (~ Ng785) ) ;
 assign n2062 = ( n426  &  Ng793 ) | ( (~ n426)  &  (~ Ng793) ) ;
 assign n2064 = ( n385  &  Ng785 ) | ( (~ n385)  &  (~ Ng785) ) ;
 assign n2066 = ( n214  &  Ng809 ) | ( (~ n214)  &  (~ Ng809) ) ;
 assign n2068 = ( n464  &  Ng801 ) | ( (~ n464)  &  (~ Ng801) ) ;
 assign n2069 = ( n279  &  Ng797 ) | ( (~ n279)  &  (~ Ng797) ) ;
 assign n2071 = ( n388  &  n627 ) | ( (~ n388)  &  (~ n627) ) ;
 assign n2072 = ( n350  &  Ng813 ) | ( (~ n350)  &  (~ Ng813) ) ;
 assign n2074 = ( n251  &  Ng789 ) | ( (~ n251)  &  (~ Ng789) ) ;
 assign n2075 = ( n464  &  n1473 ) | ( (~ n464)  &  (~ n1473) ) ;
 assign n2077 = ( (~ n385)  &  n1473 ) | ( n385  &  (~ n1473) ) ;
 assign n2078 = ( (~ n251)  &  n1473 ) | ( n251  &  (~ n1473) ) ;
 assign n2080 = ( (~ n426)  &  n1473 ) | ( n426  &  (~ n1473) ) ;
 assign n2081 = ( (~ n279)  &  n1473 ) | ( n279  &  (~ n1473) ) ;
 assign n2083 = ( n2080 ) | ( n2086 ) ;
 assign n2084 = ( n1418 ) | ( n2077 ) ;
 assign n2086 = ( n2078 ) | ( n2084 ) ;
 assign n2087 = ( n181  &  Ng105 ) | ( (~ n181)  &  (~ Ng105) ) ;
 assign n2088 = ( n298  &  Ng101 ) | ( (~ n298)  &  (~ Ng101) ) ;
 assign n2089 = ( n221  &  Ng125 ) | ( (~ n221)  &  (~ Ng125) ) ;
 assign n2090 = ( n184  &  Ng109 ) | ( (~ n184)  &  (~ Ng109) ) ;
 assign n2091 = ( n206  &  Ng121 ) | ( (~ n206)  &  (~ Ng121) ) ;
 assign n2092 = ( n195  &  Ng117 ) | ( (~ n195)  &  (~ Ng117) ) ;
 assign n2093 = ( n189  &  Ng113 ) | ( (~ n189)  &  (~ Ng113) ) ;
 assign n2094 = ( n268  &  Ng97 ) | ( (~ n268)  &  (~ Ng97) ) ;
 assign n2095 = ( n376  &  Ng105 ) | ( (~ n376)  &  (~ Ng105) ) ;
 assign n2097 = ( n335  &  Ng97 ) | ( (~ n335)  &  (~ Ng97) ) ;
 assign n2099 = ( n197  &  Ng121 ) | ( (~ n197)  &  (~ Ng121) ) ;
 assign n2101 = ( n419  &  Ng113 ) | ( (~ n419)  &  (~ Ng113) ) ;
 assign n2102 = ( n244  &  Ng109 ) | ( (~ n244)  &  (~ Ng109) ) ;
 assign n2104 = ( n338  &  n613 ) | ( (~ n338)  &  (~ n613) ) ;
 assign n2105 = ( n300  &  Ng125 ) | ( (~ n300)  &  (~ Ng125) ) ;
 assign n2107 = ( n223  &  Ng101 ) | ( (~ n223)  &  (~ Ng101) ) ;
 assign n2108 = ( n419  &  n1481 ) | ( (~ n419)  &  (~ n1481) ) ;
 assign n2110 = ( (~ n335)  &  n1481 ) | ( n335  &  (~ n1481) ) ;
 assign n2111 = ( (~ n223)  &  n1481 ) | ( n223  &  (~ n1481) ) ;
 assign n2113 = ( (~ n376)  &  n1481 ) | ( n376  &  (~ n1481) ) ;
 assign n2114 = ( (~ n244)  &  n1481 ) | ( n244  &  (~ n1481) ) ;
 assign n2116 = ( n2113 ) | ( n2119 ) ;
 assign n2117 = ( n1451 ) | ( n2110 ) ;
 assign n2119 = ( n2111 ) | ( n2117 ) ;
 assign n2121 = ( (~ n414)  &  n1339 ) | ( n414  &  (~ n1339) ) ;
 assign n2120 = ( (~ Ng2190)  &  (~ n1351) ) | ( n1349  &  (~ n1351) ) | ( (~ Ng2190)  &  n2121 ) | ( n1349  &  n2121 ) ;
 assign n2123 = ( (~ n364)  &  n1372 ) | ( n364  &  (~ n1372) ) ;
 assign n2122 = ( (~ Ng1496)  &  (~ n1384) ) | ( n1382  &  (~ n1384) ) | ( (~ Ng1496)  &  n2123 ) | ( n1382  &  n2123 ) ;
 assign n2125 = ( (~ n314)  &  n1405 ) | ( n314  &  (~ n1405) ) ;
 assign n2124 = ( (~ Ng805)  &  (~ n1417) ) | ( n1415  &  (~ n1417) ) | ( (~ Ng805)  &  n2125 ) | ( n1415  &  n2125 ) ;
 assign n2127 = ( (~ n272)  &  n1438 ) | ( n272  &  (~ n1438) ) ;
 assign n2126 = ( (~ Ng117)  &  (~ n1450) ) | ( n1448  &  (~ n1450) ) | ( (~ Ng117)  &  n2127 ) | ( n1448  &  n2127 ) ;
 assign n2138 = ( Pg3229  &  n453 ) | ( (~ Pg3229)  &  (~ n453) ) ;
 assign n2139 = ( Pg3229  &  n403 ) | ( (~ Pg3229)  &  (~ n403) ) ;
 assign n2140 = ( Pg3229  &  n353 ) | ( (~ Pg3229)  &  (~ n353) ) ;
 assign n2141 = ( Pg3229  &  n303 ) | ( (~ Pg3229)  &  (~ n303) ) ;
 assign n2143 = ( Ng13475  &  Ng2993 ) ;
 assign n2142 = ( (~ n2143)  &  Ng2998 ) | ( n2143  &  (~ Ng2998) ) ;
 assign n2145 = ( n483  &  Ng2120 ) | ( (~ n483)  &  (~ Ng2120) ) ;
 assign n2146 = ( n450  &  Ng2129 ) | ( (~ n450)  &  (~ Ng2129) ) ;
 assign n2147 = ( n295  &  Ng2124 ) | ( (~ n295)  &  (~ Ng2124) ) ;
 assign n2148 = ( n265  &  Ng2133 ) | ( (~ n265)  &  (~ Ng2133) ) ;
 assign n2149 = ( n506  &  Ng2151 ) | ( (~ n506)  &  (~ Ng2151) ) ;
 assign n2150 = ( n521  &  Ng2142 ) | ( (~ n521)  &  (~ Ng2142) ) ;
 assign n2151 = ( n414  &  Ng2138 ) | ( (~ n414)  &  (~ Ng2138) ) ;
 assign n2152 = ( n480  &  Ng2160 ) | ( (~ n480)  &  (~ Ng2160) ) ;
 assign n2153 = ( n371  &  Ng2147 ) | ( (~ n371)  &  (~ Ng2147) ) ;
 assign n2154 = ( n328  &  Ng2156 ) | ( (~ n328)  &  (~ Ng2156) ) ;
 assign n2156 = ( n438  &  Ng1426 ) | ( (~ n438)  &  (~ Ng1426) ) ;
 assign n2157 = ( n400  &  Ng1435 ) | ( (~ n400)  &  (~ Ng1435) ) ;
 assign n2158 = ( n260  &  Ng1430 ) | ( (~ n260)  &  (~ Ng1430) ) ;
 assign n2159 = ( n237  &  Ng1439 ) | ( (~ n237)  &  (~ Ng1439) ) ;
 assign n2160 = ( n471  &  Ng1457 ) | ( (~ n471)  &  (~ Ng1457) ) ;
 assign n2161 = ( n499  &  Ng1448 ) | ( (~ n499)  &  (~ Ng1448) ) ;
 assign n2162 = ( n364  &  Ng1444 ) | ( (~ n364)  &  (~ Ng1444) ) ;
 assign n2163 = ( n435  &  Ng1466 ) | ( (~ n435)  &  (~ Ng1466) ) ;
 assign n2164 = ( n321  &  Ng1453 ) | ( (~ n321)  &  (~ Ng1453) ) ;
 assign n2165 = ( n286  &  Ng1462 ) | ( (~ n286)  &  (~ Ng1462) ) ;
 assign n2167 = ( n388  &  Ng740 ) | ( (~ n388)  &  (~ Ng740) ) ;
 assign n2168 = ( n350  &  Ng749 ) | ( (~ n350)  &  (~ Ng749) ) ;
 assign n2169 = ( n232  &  Ng744 ) | ( (~ n232)  &  (~ Ng744) ) ;
 assign n2170 = ( n214  &  Ng753 ) | ( (~ n214)  &  (~ Ng753) ) ;
 assign n2171 = ( n426  &  Ng771 ) | ( (~ n426)  &  (~ Ng771) ) ;
 assign n2172 = ( n464  &  Ng762 ) | ( (~ n464)  &  (~ Ng762) ) ;
 assign n2173 = ( n314  &  Ng758 ) | ( (~ n314)  &  (~ Ng758) ) ;
 assign n2174 = ( n385  &  Ng780 ) | ( (~ n385)  &  (~ Ng780) ) ;
 assign n2175 = ( n279  &  Ng767 ) | ( (~ n279)  &  (~ Ng767) ) ;
 assign n2176 = ( n251  &  Ng776 ) | ( (~ n251)  &  (~ Ng776) ) ;
 assign n2178 = ( n338  &  Ng52 ) | ( (~ n338)  &  (~ Ng52) ) ;
 assign n2179 = ( n300  &  Ng61 ) | ( (~ n300)  &  (~ Ng61) ) ;
 assign n2180 = ( n208  &  Ng56 ) | ( (~ n208)  &  (~ Ng56) ) ;
 assign n2181 = ( n197  &  Ng65 ) | ( (~ n197)  &  (~ Ng65) ) ;
 assign n2182 = ( n376  &  Ng83 ) | ( (~ n376)  &  (~ Ng83) ) ;
 assign n2183 = ( n419  &  Ng74 ) | ( (~ n419)  &  (~ Ng74) ) ;
 assign n2184 = ( n272  &  Ng70 ) | ( (~ n272)  &  (~ Ng70) ) ;
 assign n2185 = ( n335  &  Ng92 ) | ( (~ n335)  &  (~ Ng92) ) ;
 assign n2186 = ( n244  &  Ng79 ) | ( (~ n244)  &  (~ Ng79) ) ;
 assign n2187 = ( n223  &  Ng88 ) | ( (~ n223)  &  (~ Ng88) ) ;
 assign n2189 = ( n536  &  Ng2760 ) | ( (~ n536)  &  (~ Ng2760) ) ;
 assign n2191 = ( n526  &  Ng2740 ) | ( (~ n526)  &  (~ Ng2740) ) ;
 assign n2192 = ( n532  &  Ng2753 ) | ( (~ n532)  &  (~ Ng2753) ) ;
 assign n2194 = ( n333  &  Ng2766 ) | ( (~ n333)  &  (~ Ng2766) ) ;
 assign n2196 = ( n374  &  Ng2707 ) | ( (~ n374)  &  (~ Ng2707) ) ;
 assign n2198 = ( n491  &  Ng2734 ) | ( (~ n491)  &  (~ Ng2734) ) ;
 assign n2199 = ( n417  &  Ng2727 ) | ( (~ n417)  &  (~ Ng2727) ) ;
 assign n2201 = ( n458  &  Ng2720 ) | ( (~ n458)  &  (~ Ng2720) ) ;
 assign n2203 = ( n511  &  Ng2746 ) | ( (~ n511)  &  (~ Ng2746) ) ;
 assign n2204 = ( n331  &  Ng2714 ) | ( (~ n331)  &  (~ Ng2714) ) ;
 assign n2205 = ( n528  &  Ng2066 ) | ( (~ n528)  &  (~ Ng2066) ) ;
 assign n2207 = ( n504  &  Ng2046 ) | ( (~ n504)  &  (~ Ng2046) ) ;
 assign n2208 = ( n519  &  Ng2059 ) | ( (~ n519)  &  (~ Ng2059) ) ;
 assign n2210 = ( n291  &  Ng2072 ) | ( (~ n291)  &  (~ Ng2072) ) ;
 assign n2212 = ( n324  &  Ng2013 ) | ( (~ n324)  &  (~ Ng2013) ) ;
 assign n2214 = ( n446  &  Ng2040 ) | ( (~ n446)  &  (~ Ng2040) ) ;
 assign n2215 = ( n367  &  Ng2033 ) | ( (~ n367)  &  (~ Ng2033) ) ;
 assign n2217 = ( n408  &  Ng2026 ) | ( (~ n408)  &  (~ Ng2026) ) ;
 assign n2219 = ( n476  &  Ng2052 ) | ( (~ n476)  &  (~ Ng2052) ) ;
 assign n2220 = ( n289  &  Ng2020 ) | ( (~ n289)  &  (~ Ng2020) ) ;
 assign n2221 = ( n515  &  Ng1372 ) | ( (~ n515)  &  (~ Ng1372) ) ;
 assign n2223 = ( n469  &  Ng1352 ) | ( (~ n469)  &  (~ Ng1352) ) ;
 assign n2225 = ( n497  &  Ng1365 ) | ( (~ n497)  &  (~ Ng1365) ) ;
 assign n2227 = ( n256  &  Ng1378 ) | ( (~ n256)  &  (~ Ng1378) ) ;
 assign n2229 = ( n282  &  Ng1319 ) | ( (~ n282)  &  (~ Ng1319) ) ;
 assign n2231 = ( n396  &  Ng1346 ) | ( (~ n396)  &  (~ Ng1346) ) ;
 assign n2233 = ( n317  &  Ng1339 ) | ( (~ n317)  &  (~ Ng1339) ) ;
 assign n2235 = ( n358  &  Ng1332 ) | ( (~ n358)  &  (~ Ng1332) ) ;
 assign n2237 = ( n431  &  Ng1358 ) | ( (~ n431)  &  (~ Ng1358) ) ;
 assign n2239 = ( n254  &  Ng1326 ) | ( (~ n254)  &  (~ Ng1326) ) ;
 assign n2241 = ( n493  &  Ng686 ) | ( (~ n493)  &  (~ Ng686) ) ;
 assign n2243 = ( n424  &  Ng666 ) | ( (~ n424)  &  (~ Ng666) ) ;
 assign n2245 = ( n462  &  Ng679 ) | ( (~ n462)  &  (~ Ng679) ) ;
 assign n2247 = ( n228  &  Ng692 ) | ( (~ n228)  &  (~ Ng692) ) ;
 assign n2249 = ( n247  &  Ng633 ) | ( (~ n247)  &  (~ Ng633) ) ;
 assign n2251 = ( n346  &  Ng660 ) | ( (~ n346)  &  (~ Ng660) ) ;
 assign n2253 = ( n275  &  Ng653 ) | ( (~ n275)  &  (~ Ng653) ) ;
 assign n2255 = ( n308  &  Ng646 ) | ( (~ n308)  &  (~ Ng646) ) ;
 assign n2257 = ( n381  &  Ng672 ) | ( (~ n381)  &  (~ Ng672) ) ;
 assign n2259 = ( n226  &  Ng640 ) | ( (~ n226)  &  (~ Ng640) ) ;
 assign Ng30325 = ( (~ n2730) ) ;
 assign n2278 = ( (~ n679) ) | ( n1115 ) ;
 assign Ng29445 = ( (~ n2729) ) ;
 assign n2291 = ( (~ n675) ) | ( n1091 ) ;
 assign n2295 = ( (~ n369)  &  n642 ) | ( n369  &  (~ n642) ) ;
 assign n2296 = ( (~ n412)  &  n640 ) | ( n412  &  (~ n640) ) ;
 assign n2297 = ( n1991 ) | ( n1992 ) | ( n1993 ) | ( n1988 ) | ( n1989 ) | ( n1990 ) ;
 assign n2319 = ( n1996 ) | ( n1998 ) | ( n2000 ) ;
 assign n2320 = ( n1323 ) | ( n1332 ) ;
 assign n2323 = ( (~ n1329)  &  n1330 ) ;
 assign n2324 = ( Ng2257  &  n530 ) ;
 assign n2325 = ( n414  &  n450  &  n480  &  n265  &  n521 ) ;
 assign n2326 = ( n295  &  n506  &  n2325  &  n371  &  n483  &  n328 ) ;
 assign n2327 = ( n2014 ) | ( n2015 ) ;
 assign n2330 = ( (~ n319)  &  n638 ) | ( n319  &  (~ n638) ) ;
 assign n2331 = ( (~ n362)  &  n636 ) | ( n362  &  (~ n636) ) ;
 assign n2332 = ( n2024 ) | ( n2025 ) | ( n2026 ) | ( n2021 ) | ( n2022 ) | ( n2023 ) ;
 assign n2354 = ( n2029 ) | ( n2031 ) | ( n2033 ) ;
 assign n2355 = ( n1356 ) | ( n1365 ) ;
 assign n2358 = ( (~ n1362)  &  n1363 ) ;
 assign n2359 = ( Ng2257  &  n517 ) ;
 assign n2360 = ( n364  &  n400  &  n435  &  n237  &  n499 ) ;
 assign n2361 = ( n260  &  n471  &  n2360  &  n321  &  n438  &  n286 ) ;
 assign n2362 = ( n2047 ) | ( n2048 ) ;
 assign n2365 = ( (~ n277)  &  n634 ) | ( n277  &  (~ n634) ) ;
 assign n2366 = ( (~ n312)  &  n627 ) | ( n312  &  (~ n627) ) ;
 assign n2367 = ( n2057 ) | ( n2058 ) | ( n2059 ) | ( n2054 ) | ( n2055 ) | ( n2056 ) ;
 assign n2389 = ( n2062 ) | ( n2064 ) | ( n2066 ) ;
 assign n2390 = ( n1389 ) | ( n1398 ) ;
 assign n2393 = ( (~ n1395)  &  n1396 ) ;
 assign n2394 = ( Ng2257  &  n495 ) ;
 assign n2395 = ( n314  &  n350  &  n385  &  n214  &  n464 ) ;
 assign n2396 = ( n232  &  n426  &  n2395  &  n279  &  n388  &  n251 ) ;
 assign n2397 = ( n2080 ) | ( n2081 ) ;
 assign n2400 = ( (~ n242)  &  n625 ) | ( n242  &  (~ n625) ) ;
 assign n2401 = ( (~ n270)  &  n613 ) | ( n270  &  (~ n613) ) ;
 assign n2402 = ( n2090 ) | ( n2091 ) | ( n2092 ) | ( n2087 ) | ( n2088 ) | ( n2089 ) ;
 assign n2424 = ( n2095 ) | ( n2097 ) | ( n2099 ) ;
 assign n2425 = ( n1422 ) | ( n1431 ) ;
 assign n2428 = ( (~ n1428)  &  n1429 ) ;
 assign n2429 = ( Ng2257  &  n460 ) ;
 assign n2430 = ( n272  &  n300  &  n335  &  n197  &  n419 ) ;
 assign n2431 = ( n208  &  n376  &  n2430  &  n244  &  n338  &  n223 ) ;
 assign n2432 = ( n2113 ) | ( n2114 ) ;
 assign Ng27217 = ( (~ n2728) ) ;
 assign n2444 = ( (~ n671) ) | ( n1056 ) ;
 assign n2450 = ( (~ Ng853) ) | ( (~ Ng2257) ) ;
 assign n2453 = ( Ng3139 ) | ( Ng3120 ) ;
 assign n2455 = ( Ng3126 ) | ( Ng3191 ) | ( Ng3126 ) | ( (~ Ng3110) ) ;
 assign n2460 = ( Ng3139 ) | ( (~ Ng3120) ) ;
 assign Ng23159 = ( (~ n2727) ) ;
 assign n2467 = ( (~ n667) ) | ( n1015 ) ;
 assign n2489 = ( (~ n657) ) | ( n1214 ) | ( n1540 ) ;
 assign n2491 = ( (~ n652) ) | ( n1211 ) | ( n1550 ) ;
 assign n2493 = ( (~ n647) ) | ( n1208 ) | ( n1560 ) ;
 assign n2495 = ( (~ n645) ) | ( n1205 ) | ( n1570 ) ;
 assign n2497 = ( n2453 ) | ( n1768 ) | ( Ng3135 ) | ( Ng3147 ) ;
 assign n2498 = ( Ng3147 ) | ( n2455 ) ;
 assign n2499 = ( (~ Ng3139) ) | ( Ng3120 ) ;
 assign n2500 = ( (~ Ng3135) ) | ( n2498 ) ;
 assign n2501 = ( n2499 ) | ( n2500 ) ;
 assign n2502 = ( n1524 ) | ( n2498 ) ;
 assign n2503 = ( (~ Ng3139) ) | ( (~ Ng3120) ) ;
 assign n2504 = ( n2500 ) | ( n2503 ) ;
 assign n2505 = ( Ng3135 ) | ( n2498 ) ;
 assign n2506 = ( n2453 ) | ( n2505 ) ;
 assign n2508 = ( n2499 ) | ( n2505 ) ;
 assign n2510 = ( n2460 ) | ( n2505 ) ;
 assign n2512 = ( n2503 ) | ( n2505 ) ;
 assign n2514 = ( (~ Ng3147) ) | ( n2455 ) | ( Ng3135 ) ;
 assign n2515 = ( n2453 ) | ( n2514 ) ;
 assign n2517 = ( n2499 ) | ( n2514 ) ;
 assign n2519 = ( n2460 ) | ( n2514 ) ;
 assign n2520 = ( n2503 ) | ( n2514 ) ;
 assign n2521 = ( n2453 ) | ( n2500 ) ;
 assign n2523 = ( Ng2740  &  Ng2746  &  n1871 ) ;
 assign n2524 = ( Ng2998  &  Ng3024  &  Ng3013  &  Ng3002  &  (~ Ng2993)  &  (~ Ng3006)  &  (~ Ng3010) ) ;
 assign n2534 = ( (~ n611) ) | ( (~ n632) ) ;
 assign n2546 = ( n109  &  (~ n611)  &  (~ n1630) ) ;
 assign n2545 = ( n2546 ) | ( n1639 ) | ( n1641 ) ;
 assign n2547 = ( (~ Ng3032)  &  Ng3018  &  (~ Ng3036)  &  n2524  &  Ng3028 ) ;
 assign n2551 = ( Ng2046  &  Ng2052  &  n1875 ) ;
 assign n2560 = ( (~ n597) ) | ( (~ n618) ) ;
 assign n2572 = ( n100  &  (~ n597)  &  (~ n1665) ) ;
 assign n2571 = ( n2572 ) | ( n1674 ) | ( n1676 ) ;
 assign n2575 = ( Ng1352  &  Ng1358  &  n1879 ) ;
 assign n2584 = ( (~ n583) ) | ( (~ n604) ) ;
 assign n2596 = ( n88  &  (~ n583)  &  (~ n1700) ) ;
 assign n2595 = ( n2596 ) | ( n1709 ) | ( n1711 ) ;
 assign n2599 = ( Ng666  &  Ng672  &  n1883 ) ;
 assign n2608 = ( (~ n574) ) | ( (~ n590) ) ;
 assign n2620 = ( n76  &  (~ n574)  &  (~ n1735) ) ;
 assign n2619 = ( n2620 ) | ( n1744 ) | ( n1746 ) ;
 assign n2653 = ( n455  &  n4136 ) | ( (~ n488)  &  n4136 ) | ( (~ n1786)  &  n4136 ) ;
 assign n2662 = ( n405  &  n4137 ) | ( (~ n443)  &  n4137 ) | ( (~ n1797)  &  n4137 ) ;
 assign n2671 = ( n355  &  n4138 ) | ( (~ n393)  &  n4138 ) | ( (~ n1807)  &  n4138 ) ;
 assign n2680 = ( n305  &  n4139 ) | ( (~ n343)  &  n4139 ) | ( (~ n1817)  &  n4139 ) ;
 assign n2694 = ( Ng2998  &  n2143 ) ;
 assign n2695 = ( (~ Ng3002) ) | ( (~ n2694) ) | ( (~ Ng3006) ) ;
 assign n2699 = ( Ng2892  &  Ng2896  &  n1934 ) ;
 assign n2702 = ( Ng2599  &  (~ Ng2733)  &  Ng2612 ) ;
 assign n2703 = ( n721 ) | ( Ng2912 ) | ( Ng2920 ) | ( (~ Ng2924) ) | ( (~ Ng2883) ) | ( Ng2888 ) | ( Ng2917 ) ;
 assign n2704 = ( Ng1905  &  (~ Ng2039)  &  Ng1918 ) ;
 assign n2705 = ( Ng1211  &  (~ Ng1345)  &  Ng1224 ) ;
 assign n2706 = ( Ng525  &  (~ Ng659)  &  Ng538 ) ;
 assign n2710 = ( (~ n480)  &  n1352 ) | ( n480  &  (~ n1352) ) ;
 assign n2711 = ( (~ n435)  &  n1385 ) | ( n435  &  (~ n1385) ) ;
 assign n2712 = ( (~ n385)  &  n1418 ) | ( n385  &  (~ n1418) ) ;
 assign n2713 = ( (~ n335)  &  n1451 ) | ( n335  &  (~ n1451) ) ;
 assign n2714 = ( (~ Ng3024)  &  n1865 ) | ( Ng3024  &  (~ n1865) ) ;
 assign n2715 = ( (~ n455)  &  n1786 ) | ( n455  &  (~ n1786) ) ;
 assign n2716 = ( (~ n405)  &  n1797 ) | ( n405  &  (~ n1797) ) ;
 assign n2717 = ( (~ n355)  &  n1807 ) | ( n355  &  (~ n1807) ) ;
 assign n2718 = ( (~ n305)  &  n1817 ) | ( n305  &  (~ n1817) ) ;
 assign n2721 = ( (~ n1137)  &  n1146 ) | ( n1137  &  (~ n1146) ) ;
 assign Ng21966 = ( (~ Ng3083)  &  n2721 ) | ( Ng3083  &  (~ n2721) ) ;
 assign n2722 = ( (~ n1140)  &  n1143 ) | ( n1140  &  (~ n1143) ) ;
 assign Ng21964 = ( (~ Ng2990)  &  n2722 ) | ( Ng2990  &  (~ n2722) ) ;
 assign Ng20604 = ( n2721  &  n4898 ) | ( (~ n2721)  &  (~ n4898) ) ;
 assign Ng20594 = ( n2722  &  n4898 ) | ( (~ n2722)  &  (~ n4898) ) ;
 assign n2724 = ( (~ n1127)  &  n1132 ) | ( n1127  &  (~ n1132) ) ;
 assign Ng19061 = ( (~ Ng2934)  &  n2724 ) | ( Ng2934  &  (~ n2724) ) ;
 assign n2725 = ( (~ n1117)  &  n1122 ) | ( n1117  &  (~ n1122) ) ;
 assign Ng19060 = ( (~ Ng2962)  &  n2725 ) | ( Ng2962  &  (~ n2725) ) ;
 assign n2726 = ( n536  &  (~ n569) ) | ( (~ n536)  &  (~ n3742) ) | ( (~ n569)  &  (~ n3742) ) ;
 assign n2727 = ( (~ Ng8284)  &  n3884 ) | ( (~ Ng544)  &  n3884 ) ;
 assign n2728 = ( (~ Ng8293)  &  n3886 ) | ( Ng8293  &  (~ Ng1230) ) | ( n3886  &  (~ Ng1230) ) ;
 assign n2729 = ( (~ Ng8302)  &  n3889 ) | ( Ng8302  &  (~ Ng1924) ) | ( n3889  &  (~ Ng1924) ) ;
 assign n2730 = ( (~ Ng8311)  &  n3892 ) | ( Ng8311  &  (~ Ng2618) ) | ( n3892  &  (~ Ng2618) ) ;
 assign n2731 = ( n333  &  (~ n662) ) | ( (~ n333)  &  n3743 ) | ( (~ n662)  &  n3743 ) ;
 assign n2732 = ( n374  &  (~ n662) ) | ( (~ n374)  &  n3743 ) | ( (~ n662)  &  n3743 ) ;
 assign n2733 = ( n458  &  (~ n662) ) | ( (~ n458)  &  n3743 ) | ( (~ n662)  &  n3743 ) ;
 assign n2734 = ( n417  &  (~ n569) ) | ( (~ n417)  &  (~ n3742) ) | ( (~ n569)  &  (~ n3742) ) ;
 assign n2735 = ( (~ Ng1315)  &  (~ Ng3108) ) | ( Ng1315  &  n2730 ) | ( (~ Ng3108)  &  n2730 ) ;
 assign Ng30943 = ( (~ n2735) ) ;
 assign n2736 = ( (~ wire1603)  &  (~ Ng3107) ) | ( wire1603  &  n2730 ) | ( (~ Ng3107)  &  n2730 ) ;
 assign Ng30942 = ( (~ n2736) ) ;
 assign n2737 = ( (~ wire1605)  &  (~ Ng3106) ) | ( wire1605  &  n2730 ) | ( (~ Ng3106)  &  n2730 ) ;
 assign Ng30941 = ( (~ n2737) ) ;
 assign n2738 = ( n528  &  (~ n564) ) | ( (~ n528)  &  (~ n3740) ) | ( (~ n564)  &  (~ n3740) ) ;
 assign n2739 = ( n291  &  (~ n659) ) | ( (~ n291)  &  n3741 ) | ( (~ n659)  &  n3741 ) ;
 assign n2740 = ( n324  &  (~ n659) ) | ( (~ n324)  &  n3741 ) | ( (~ n659)  &  n3741 ) ;
 assign n2741 = ( n408  &  (~ n659) ) | ( (~ n408)  &  n3741 ) | ( (~ n659)  &  n3741 ) ;
 assign n2742 = ( n367  &  (~ n564) ) | ( (~ n367)  &  (~ n3740) ) | ( (~ n564)  &  (~ n3740) ) ;
 assign n2743 = ( (~ Ng853)  &  (~ Ng2392) ) | ( Ng853  &  n3916 ) | ( (~ Ng2392)  &  n3916 ) ;
 assign Ng30907 = ( (~ n2743) ) ;
 assign n2744 = ( (~ wire1594)  &  (~ Ng2391) ) | ( wire1594  &  n3916 ) | ( (~ Ng2391)  &  n3916 ) ;
 assign Ng30906 = ( (~ n2744) ) ;
 assign n2745 = ( (~ wire1612)  &  (~ Ng2390) ) | ( wire1612  &  n3916 ) | ( (~ Ng2390)  &  n3916 ) ;
 assign Ng30905 = ( (~ n2745) ) ;
 assign n2746 = ( (~ n295)  &  (~ n328)  &  (~ n371)  &  (~ n483)  &  (~ n506)  &  n2325 ) ;
 assign n2747 = ( n1457  &  n2326 ) | ( (~ n1457)  &  n2746 ) | ( n2326  &  n2746 ) ;
 assign n2748 = ( Ng853  &  (~ n986) ) | ( (~ Ng853)  &  (~ Ng2348) ) | ( (~ n986)  &  (~ Ng2348) ) ;
 assign Ng30904 = ( (~ n2748) ) ;
 assign n2749 = ( wire1594  &  (~ n986) ) | ( (~ wire1594)  &  (~ Ng2345) ) | ( (~ n986)  &  (~ Ng2345) ) ;
 assign Ng30903 = ( (~ n2749) ) ;
 assign n2750 = ( wire1612  &  (~ n986) ) | ( (~ wire1612)  &  (~ Ng2342) ) | ( (~ n986)  &  (~ Ng2342) ) ;
 assign Ng30902 = ( (~ n2750) ) ;
 assign n2751 = ( Ng853  &  (~ n968) ) | ( (~ Ng853)  &  (~ Ng2321) ) | ( (~ n968)  &  (~ Ng2321) ) ;
 assign Ng30901 = ( (~ n2751) ) ;
 assign n2752 = ( wire1594  &  (~ n968) ) | ( (~ wire1594)  &  (~ Ng2318) ) | ( (~ n968)  &  (~ Ng2318) ) ;
 assign Ng30900 = ( (~ n2752) ) ;
 assign n2753 = ( wire1612  &  (~ n968) ) | ( (~ wire1612)  &  (~ Ng2315) ) | ( (~ n968)  &  (~ Ng2315) ) ;
 assign Ng30899 = ( (~ n2753) ) ;
 assign n2754 = ( Ng853  &  (~ n962) ) | ( (~ Ng853)  &  (~ Ng2312) ) | ( (~ n962)  &  (~ Ng2312) ) ;
 assign Ng30898 = ( (~ n2754) ) ;
 assign n2755 = ( wire1594  &  (~ n962) ) | ( (~ wire1594)  &  (~ Ng2309) ) | ( (~ n962)  &  (~ Ng2309) ) ;
 assign Ng30897 = ( (~ n2755) ) ;
 assign n2756 = ( wire1612  &  (~ n962) ) | ( (~ wire1612)  &  (~ Ng2306) ) | ( (~ n962)  &  (~ Ng2306) ) ;
 assign Ng30896 = ( (~ n2756) ) ;
 assign n2757 = ( Ng853  &  (~ n954) ) | ( (~ Ng853)  &  (~ Ng2303) ) | ( (~ n954)  &  (~ Ng2303) ) ;
 assign Ng30895 = ( (~ n2757) ) ;
 assign n2758 = ( wire1594  &  (~ n954) ) | ( (~ wire1594)  &  (~ Ng2300) ) | ( (~ n954)  &  (~ Ng2300) ) ;
 assign Ng30894 = ( (~ n2758) ) ;
 assign n2759 = ( wire1612  &  (~ n954) ) | ( (~ wire1612)  &  (~ Ng2297) ) | ( (~ n954)  &  (~ Ng2297) ) ;
 assign Ng30893 = ( (~ n2759) ) ;
 assign n2760 = ( Ng853  &  (~ n989) ) | ( (~ Ng853)  &  (~ Ng2276) ) | ( (~ n989)  &  (~ Ng2276) ) ;
 assign Ng30892 = ( (~ n2760) ) ;
 assign n2761 = ( wire1594  &  (~ n989) ) | ( (~ wire1594)  &  (~ Ng2273) ) | ( (~ n989)  &  (~ Ng2273) ) ;
 assign Ng30891 = ( (~ n2761) ) ;
 assign n2762 = ( wire1612  &  (~ n989) ) | ( (~ wire1612)  &  (~ Ng2270) ) | ( (~ n989)  &  (~ Ng2270) ) ;
 assign Ng30890 = ( (~ n2762) ) ;
 assign n2763 = ( (~ Ng853)  &  (~ Ng1698) ) | ( Ng853  &  n3932 ) | ( (~ Ng1698)  &  n3932 ) ;
 assign Ng30889 = ( (~ n2763) ) ;
 assign n2764 = ( (~ wire1594)  &  (~ Ng1697) ) | ( wire1594  &  n3932 ) | ( (~ Ng1697)  &  n3932 ) ;
 assign Ng30888 = ( (~ n2764) ) ;
 assign n2765 = ( (~ wire1612)  &  (~ Ng1696) ) | ( wire1612  &  n3932 ) | ( (~ Ng1696)  &  n3932 ) ;
 assign Ng30887 = ( (~ n2765) ) ;
 assign n2766 = ( (~ n260)  &  (~ n286)  &  (~ n321)  &  (~ n438)  &  (~ n471)  &  n2360 ) ;
 assign n2767 = ( n1465  &  n2361 ) | ( (~ n1465)  &  n2766 ) | ( n2361  &  n2766 ) ;
 assign n2768 = ( Ng853  &  (~ n980) ) | ( (~ Ng853)  &  (~ Ng1654) ) | ( (~ n980)  &  (~ Ng1654) ) ;
 assign Ng30886 = ( (~ n2768) ) ;
 assign n2769 = ( wire1594  &  (~ n980) ) | ( (~ wire1594)  &  (~ Ng1651) ) | ( (~ n980)  &  (~ Ng1651) ) ;
 assign Ng30885 = ( (~ n2769) ) ;
 assign n2770 = ( wire1612  &  (~ n980) ) | ( (~ wire1612)  &  (~ Ng1648) ) | ( (~ n980)  &  (~ Ng1648) ) ;
 assign Ng30884 = ( (~ n2770) ) ;
 assign n2771 = ( Ng853  &  (~ n959) ) | ( (~ Ng853)  &  (~ Ng1627) ) | ( (~ n959)  &  (~ Ng1627) ) ;
 assign Ng30883 = ( (~ n2771) ) ;
 assign n2772 = ( wire1594  &  (~ n959) ) | ( (~ wire1594)  &  (~ Ng1624) ) | ( (~ n959)  &  (~ Ng1624) ) ;
 assign Ng30882 = ( (~ n2772) ) ;
 assign n2773 = ( wire1612  &  (~ n959) ) | ( (~ wire1612)  &  (~ Ng1621) ) | ( (~ n959)  &  (~ Ng1621) ) ;
 assign Ng30881 = ( (~ n2773) ) ;
 assign n2774 = ( Ng853  &  (~ n951) ) | ( (~ Ng853)  &  (~ Ng1618) ) | ( (~ n951)  &  (~ Ng1618) ) ;
 assign Ng30880 = ( (~ n2774) ) ;
 assign n2775 = ( wire1594  &  (~ n951) ) | ( (~ wire1594)  &  (~ Ng1615) ) | ( (~ n951)  &  (~ Ng1615) ) ;
 assign Ng30879 = ( (~ n2775) ) ;
 assign n2776 = ( wire1612  &  (~ n951) ) | ( (~ wire1612)  &  (~ Ng1612) ) | ( (~ n951)  &  (~ Ng1612) ) ;
 assign Ng30878 = ( (~ n2776) ) ;
 assign n2777 = ( Ng853  &  (~ n943) ) | ( (~ Ng853)  &  (~ Ng1609) ) | ( (~ n943)  &  (~ Ng1609) ) ;
 assign Ng30877 = ( (~ n2777) ) ;
 assign n2778 = ( wire1594  &  (~ n943) ) | ( (~ wire1594)  &  (~ Ng1606) ) | ( (~ n943)  &  (~ Ng1606) ) ;
 assign Ng30876 = ( (~ n2778) ) ;
 assign n2779 = ( wire1612  &  (~ n943) ) | ( (~ wire1612)  &  (~ Ng1603) ) | ( (~ n943)  &  (~ Ng1603) ) ;
 assign Ng30875 = ( (~ n2779) ) ;
 assign n2780 = ( Ng853  &  (~ n983) ) | ( (~ Ng853)  &  (~ Ng1582) ) | ( (~ n983)  &  (~ Ng1582) ) ;
 assign Ng30874 = ( (~ n2780) ) ;
 assign n2781 = ( wire1594  &  (~ n983) ) | ( (~ wire1594)  &  (~ Ng1579) ) | ( (~ n983)  &  (~ Ng1579) ) ;
 assign Ng30873 = ( (~ n2781) ) ;
 assign n2782 = ( wire1612  &  (~ n983) ) | ( (~ wire1612)  &  (~ Ng1576) ) | ( (~ n983)  &  (~ Ng1576) ) ;
 assign Ng30872 = ( (~ n2782) ) ;
 assign n2783 = ( (~ Ng853)  &  (~ Ng1004) ) | ( Ng853  &  n3948 ) | ( (~ Ng1004)  &  n3948 ) ;
 assign Ng30871 = ( (~ n2783) ) ;
 assign n2784 = ( (~ wire1594)  &  (~ Ng1003) ) | ( wire1594  &  n3948 ) | ( (~ Ng1003)  &  n3948 ) ;
 assign Ng30870 = ( (~ n2784) ) ;
 assign n2785 = ( (~ wire1612)  &  (~ Ng1002) ) | ( wire1612  &  n3948 ) | ( (~ Ng1002)  &  n3948 ) ;
 assign Ng30869 = ( (~ n2785) ) ;
 assign n2786 = ( (~ n232)  &  (~ n251)  &  (~ n279)  &  (~ n388)  &  (~ n426)  &  n2395 ) ;
 assign n2787 = ( n1473  &  n2396 ) | ( (~ n1473)  &  n2786 ) | ( n2396  &  n2786 ) ;
 assign n2788 = ( Ng853  &  (~ n974) ) | ( (~ Ng853)  &  (~ Ng960) ) | ( (~ n974)  &  (~ Ng960) ) ;
 assign Ng30868 = ( (~ n2788) ) ;
 assign n2789 = ( wire1594  &  (~ n974) ) | ( (~ wire1594)  &  (~ Ng957) ) | ( (~ n974)  &  (~ Ng957) ) ;
 assign Ng30867 = ( (~ n2789) ) ;
 assign n2790 = ( wire1612  &  (~ n974) ) | ( (~ wire1612)  &  (~ Ng954) ) | ( (~ n974)  &  (~ Ng954) ) ;
 assign Ng30866 = ( (~ n2790) ) ;
 assign n2791 = ( Ng853  &  (~ n948) ) | ( (~ Ng853)  &  (~ Ng933) ) | ( (~ n948)  &  (~ Ng933) ) ;
 assign Ng30865 = ( (~ n2791) ) ;
 assign n2792 = ( wire1594  &  (~ n948) ) | ( (~ wire1594)  &  (~ Ng930) ) | ( (~ n948)  &  (~ Ng930) ) ;
 assign Ng30864 = ( (~ n2792) ) ;
 assign n2793 = ( wire1612  &  (~ n948) ) | ( (~ wire1612)  &  (~ Ng927) ) | ( (~ n948)  &  (~ Ng927) ) ;
 assign Ng30863 = ( (~ n2793) ) ;
 assign n2794 = ( Ng853  &  (~ n940) ) | ( (~ Ng853)  &  (~ Ng924) ) | ( (~ n940)  &  (~ Ng924) ) ;
 assign Ng30862 = ( (~ n2794) ) ;
 assign n2795 = ( wire1594  &  (~ n940) ) | ( (~ wire1594)  &  (~ Ng921) ) | ( (~ n940)  &  (~ Ng921) ) ;
 assign Ng30861 = ( (~ n2795) ) ;
 assign n2796 = ( wire1612  &  (~ n940) ) | ( (~ wire1612)  &  (~ Ng918) ) | ( (~ n940)  &  (~ Ng918) ) ;
 assign Ng30860 = ( (~ n2796) ) ;
 assign n2797 = ( Ng853  &  (~ n932) ) | ( (~ Ng853)  &  (~ Ng915) ) | ( (~ n932)  &  (~ Ng915) ) ;
 assign Ng30859 = ( (~ n2797) ) ;
 assign n2798 = ( wire1594  &  (~ n932) ) | ( (~ wire1594)  &  (~ Ng912) ) | ( (~ n932)  &  (~ Ng912) ) ;
 assign Ng30858 = ( (~ n2798) ) ;
 assign n2799 = ( wire1612  &  (~ n932) ) | ( (~ wire1612)  &  (~ Ng909) ) | ( (~ n932)  &  (~ Ng909) ) ;
 assign Ng30857 = ( (~ n2799) ) ;
 assign n2800 = ( Ng853  &  (~ n977) ) | ( (~ Ng853)  &  (~ Ng888) ) | ( (~ n977)  &  (~ Ng888) ) ;
 assign Ng30856 = ( (~ n2800) ) ;
 assign n2801 = ( wire1594  &  (~ n977) ) | ( (~ wire1594)  &  (~ Ng885) ) | ( (~ n977)  &  (~ Ng885) ) ;
 assign Ng30855 = ( (~ n2801) ) ;
 assign n2802 = ( wire1612  &  (~ n977) ) | ( (~ wire1612)  &  (~ Ng882) ) | ( (~ n977)  &  (~ Ng882) ) ;
 assign Ng30854 = ( (~ n2802) ) ;
 assign n2803 = ( (~ Ng853)  &  (~ Ng317) ) | ( Ng853  &  n3964 ) | ( (~ Ng317)  &  n3964 ) ;
 assign Ng30853 = ( (~ n2803) ) ;
 assign n2804 = ( (~ wire1594)  &  (~ Ng316) ) | ( wire1594  &  n3964 ) | ( (~ Ng316)  &  n3964 ) ;
 assign Ng30852 = ( (~ n2804) ) ;
 assign n2805 = ( (~ wire1612)  &  (~ Ng315) ) | ( wire1612  &  n3964 ) | ( (~ Ng315)  &  n3964 ) ;
 assign Ng30851 = ( (~ n2805) ) ;
 assign n2806 = ( (~ n208)  &  (~ n223)  &  (~ n244)  &  (~ n338)  &  (~ n376)  &  n2430 ) ;
 assign n2807 = ( n1481  &  n2431 ) | ( (~ n1481)  &  n2806 ) | ( n2431  &  n2806 ) ;
 assign n2808 = ( Ng853  &  (~ n965) ) | ( (~ Ng853)  &  (~ Ng273) ) | ( (~ n965)  &  (~ Ng273) ) ;
 assign Ng30850 = ( (~ n2808) ) ;
 assign n2809 = ( wire1594  &  (~ n965) ) | ( (~ wire1594)  &  (~ Ng270) ) | ( (~ n965)  &  (~ Ng270) ) ;
 assign Ng30849 = ( (~ n2809) ) ;
 assign n2810 = ( wire1612  &  (~ n965) ) | ( (~ wire1612)  &  (~ Ng267) ) | ( (~ n965)  &  (~ Ng267) ) ;
 assign Ng30848 = ( (~ n2810) ) ;
 assign n2811 = ( Ng853  &  (~ n937) ) | ( (~ Ng853)  &  (~ Ng246) ) | ( (~ n937)  &  (~ Ng246) ) ;
 assign Ng30847 = ( (~ n2811) ) ;
 assign n2812 = ( wire1594  &  (~ n937) ) | ( (~ wire1594)  &  (~ Ng243) ) | ( (~ n937)  &  (~ Ng243) ) ;
 assign Ng30846 = ( (~ n2812) ) ;
 assign n2813 = ( wire1612  &  (~ n937) ) | ( (~ wire1612)  &  (~ Ng240) ) | ( (~ n937)  &  (~ Ng240) ) ;
 assign Ng30845 = ( (~ n2813) ) ;
 assign n2814 = ( Ng853  &  (~ n929) ) | ( (~ Ng853)  &  (~ Ng237) ) | ( (~ n929)  &  (~ Ng237) ) ;
 assign Ng30844 = ( (~ n2814) ) ;
 assign n2815 = ( wire1594  &  (~ n929) ) | ( (~ wire1594)  &  (~ Ng234) ) | ( (~ n929)  &  (~ Ng234) ) ;
 assign Ng30843 = ( (~ n2815) ) ;
 assign n2816 = ( wire1612  &  (~ n929) ) | ( (~ wire1612)  &  (~ Ng231) ) | ( (~ n929)  &  (~ Ng231) ) ;
 assign Ng30842 = ( (~ n2816) ) ;
 assign n2817 = ( Ng853  &  (~ n924) ) | ( (~ Ng853)  &  (~ Ng228) ) | ( (~ n924)  &  (~ Ng228) ) ;
 assign Ng30841 = ( (~ n2817) ) ;
 assign n2818 = ( wire1594  &  (~ n924) ) | ( (~ wire1594)  &  (~ Ng225) ) | ( (~ n924)  &  (~ Ng225) ) ;
 assign Ng30840 = ( (~ n2818) ) ;
 assign n2819 = ( wire1612  &  (~ n924) ) | ( (~ wire1612)  &  (~ Ng222) ) | ( (~ n924)  &  (~ Ng222) ) ;
 assign Ng30839 = ( (~ n2819) ) ;
 assign n2820 = ( Ng853  &  (~ n971) ) | ( (~ Ng853)  &  (~ Ng201) ) | ( (~ n971)  &  (~ Ng201) ) ;
 assign Ng30838 = ( (~ n2820) ) ;
 assign n2821 = ( wire1594  &  (~ n971) ) | ( (~ wire1594)  &  (~ Ng198) ) | ( (~ n971)  &  (~ Ng198) ) ;
 assign Ng30837 = ( (~ n2821) ) ;
 assign n2822 = ( wire1612  &  (~ n971) ) | ( (~ wire1612)  &  (~ Ng195) ) | ( (~ n971)  &  (~ Ng195) ) ;
 assign Ng30836 = ( (~ n2822) ) ;
 assign n2823 = ( Ng853  &  (~ n919) ) | ( (~ Ng853)  &  (~ Ng2395) ) | ( (~ n919)  &  (~ Ng2395) ) ;
 assign Ng30721 = ( (~ n2823) ) ;
 assign n2824 = ( (~ wire1594)  &  (~ Ng2394) ) | ( wire1594  &  (~ n919) ) | ( (~ Ng2394)  &  (~ n919) ) ;
 assign Ng30720 = ( (~ n2824) ) ;
 assign n2825 = ( wire1612  &  (~ n919) ) | ( (~ wire1612)  &  (~ Ng2393) ) | ( (~ n919)  &  (~ Ng2393) ) ;
 assign Ng30719 = ( (~ n2825) ) ;
 assign n2826 = ( Ng853  &  (~ n914) ) | ( (~ Ng853)  &  (~ Ng1701) ) | ( (~ n914)  &  (~ Ng1701) ) ;
 assign Ng30718 = ( (~ n2826) ) ;
 assign n2827 = ( (~ wire1594)  &  (~ Ng1700) ) | ( wire1594  &  (~ n914) ) | ( (~ Ng1700)  &  (~ n914) ) ;
 assign Ng30717 = ( (~ n2827) ) ;
 assign n2828 = ( wire1612  &  (~ n914) ) | ( (~ wire1612)  &  (~ Ng1699) ) | ( (~ n914)  &  (~ Ng1699) ) ;
 assign Ng30716 = ( (~ n2828) ) ;
 assign n2829 = ( Ng853  &  (~ n909) ) | ( (~ Ng853)  &  (~ Ng1007) ) | ( (~ n909)  &  (~ Ng1007) ) ;
 assign Ng30715 = ( (~ n2829) ) ;
 assign n2830 = ( (~ wire1594)  &  (~ Ng1006) ) | ( wire1594  &  (~ n909) ) | ( (~ Ng1006)  &  (~ n909) ) ;
 assign Ng30714 = ( (~ n2830) ) ;
 assign n2831 = ( wire1612  &  (~ n909) ) | ( (~ wire1612)  &  (~ Ng1005) ) | ( (~ n909)  &  (~ Ng1005) ) ;
 assign Ng30713 = ( (~ n2831) ) ;
 assign n2832 = ( Ng853  &  (~ n904) ) | ( (~ Ng853)  &  (~ Ng320) ) | ( (~ n904)  &  (~ Ng320) ) ;
 assign Ng30712 = ( (~ n2832) ) ;
 assign n2833 = ( (~ wire1594)  &  (~ Ng319) ) | ( wire1594  &  (~ n904) ) | ( (~ Ng319)  &  (~ n904) ) ;
 assign Ng30711 = ( (~ n2833) ) ;
 assign n2834 = ( wire1612  &  (~ n904) ) | ( (~ wire1612)  &  (~ Ng318) ) | ( (~ n904)  &  (~ Ng318) ) ;
 assign Ng30710 = ( (~ n2834) ) ;
 assign n2836 = ( (~ n1351)  &  n1459 ) | ( n1351  &  n3993 ) | ( n1459  &  n3993 ) ;
 assign n2837 = ( (~ Ng853)  &  (~ Ng2339) ) | ( Ng853  &  (~ n2836) ) | ( (~ Ng2339)  &  (~ n2836) ) ;
 assign Ng30565 = ( (~ n2837) ) ;
 assign n2838 = ( (~ wire1594)  &  (~ Ng2336) ) | ( wire1594  &  (~ n2836) ) | ( (~ Ng2336)  &  (~ n2836) ) ;
 assign Ng30564 = ( (~ n2838) ) ;
 assign n2839 = ( (~ wire1612)  &  (~ Ng2333) ) | ( wire1612  &  (~ n2836) ) | ( (~ Ng2333)  &  (~ n2836) ) ;
 assign Ng30563 = ( (~ n2839) ) ;
 assign n2840 = ( Ng853  &  n2120 ) | ( (~ Ng853)  &  (~ Ng2330) ) | ( n2120  &  (~ Ng2330) ) ;
 assign Ng30562 = ( (~ n2840) ) ;
 assign n2841 = ( wire1594  &  n2120 ) | ( (~ wire1594)  &  (~ Ng2327) ) | ( n2120  &  (~ Ng2327) ) ;
 assign Ng30561 = ( (~ n2841) ) ;
 assign n2842 = ( wire1612  &  n2120 ) | ( (~ wire1612)  &  (~ Ng2324) ) | ( n2120  &  (~ Ng2324) ) ;
 assign Ng30560 = ( (~ n2842) ) ;
 assign n2844 = ( (~ n1351)  &  n1460 ) | ( n1351  &  n3994 ) | ( n1460  &  n3994 ) ;
 assign n2845 = ( (~ Ng853)  &  (~ Ng2294) ) | ( Ng853  &  (~ n2844) ) | ( (~ Ng2294)  &  (~ n2844) ) ;
 assign Ng30559 = ( (~ n2845) ) ;
 assign n2846 = ( (~ wire1594)  &  (~ Ng2291) ) | ( wire1594  &  (~ n2844) ) | ( (~ Ng2291)  &  (~ n2844) ) ;
 assign Ng30558 = ( (~ n2846) ) ;
 assign n2847 = ( (~ wire1612)  &  (~ Ng2288) ) | ( wire1612  &  (~ n2844) ) | ( (~ Ng2288)  &  (~ n2844) ) ;
 assign Ng30557 = ( (~ n2847) ) ;
 assign n2849 = ( (~ n1351)  &  n1461 ) | ( n1351  &  n3995 ) | ( n1461  &  n3995 ) ;
 assign n2850 = ( (~ Ng853)  &  (~ Ng2285) ) | ( Ng853  &  (~ n2849) ) | ( (~ Ng2285)  &  (~ n2849) ) ;
 assign Ng30556 = ( (~ n2850) ) ;
 assign n2851 = ( (~ wire1594)  &  (~ Ng2282) ) | ( wire1594  &  (~ n2849) ) | ( (~ Ng2282)  &  (~ n2849) ) ;
 assign Ng30555 = ( (~ n2851) ) ;
 assign n2852 = ( (~ wire1612)  &  (~ Ng2279) ) | ( wire1612  &  (~ n2849) ) | ( (~ Ng2279)  &  (~ n2849) ) ;
 assign Ng30554 = ( (~ n2852) ) ;
 assign n2854 = ( (~ n1351)  &  n1462 ) | ( n1351  &  n2710 ) | ( n1462  &  n2710 ) ;
 assign n2855 = ( (~ Ng853)  &  (~ Ng2267) ) | ( Ng853  &  (~ n2854) ) | ( (~ Ng2267)  &  (~ n2854) ) ;
 assign Ng30553 = ( (~ n2855) ) ;
 assign n2856 = ( (~ wire1594)  &  (~ Ng2264) ) | ( wire1594  &  (~ n2854) ) | ( (~ Ng2264)  &  (~ n2854) ) ;
 assign Ng30552 = ( (~ n2856) ) ;
 assign n2857 = ( (~ wire1612)  &  (~ Ng2261) ) | ( wire1612  &  (~ n2854) ) | ( (~ Ng2261)  &  (~ n2854) ) ;
 assign Ng30551 = ( (~ n2857) ) ;
 assign n2859 = ( (~ n1384)  &  n1467 ) | ( n1384  &  n3997 ) | ( n1467  &  n3997 ) ;
 assign n2860 = ( (~ Ng853)  &  (~ Ng1645) ) | ( Ng853  &  (~ n2859) ) | ( (~ Ng1645)  &  (~ n2859) ) ;
 assign Ng30550 = ( (~ n2860) ) ;
 assign n2861 = ( (~ wire1594)  &  (~ Ng1642) ) | ( wire1594  &  (~ n2859) ) | ( (~ Ng1642)  &  (~ n2859) ) ;
 assign Ng30549 = ( (~ n2861) ) ;
 assign n2862 = ( (~ wire1612)  &  (~ Ng1639) ) | ( wire1612  &  (~ n2859) ) | ( (~ Ng1639)  &  (~ n2859) ) ;
 assign Ng30548 = ( (~ n2862) ) ;
 assign n2863 = ( Ng853  &  n2122 ) | ( (~ Ng853)  &  (~ Ng1636) ) | ( n2122  &  (~ Ng1636) ) ;
 assign Ng30547 = ( (~ n2863) ) ;
 assign n2864 = ( wire1594  &  n2122 ) | ( (~ wire1594)  &  (~ Ng1633) ) | ( n2122  &  (~ Ng1633) ) ;
 assign Ng30546 = ( (~ n2864) ) ;
 assign n2865 = ( wire1612  &  n2122 ) | ( (~ wire1612)  &  (~ Ng1630) ) | ( n2122  &  (~ Ng1630) ) ;
 assign Ng30545 = ( (~ n2865) ) ;
 assign n2867 = ( (~ n1384)  &  n1468 ) | ( n1384  &  n3998 ) | ( n1468  &  n3998 ) ;
 assign n2868 = ( (~ Ng853)  &  (~ Ng1600) ) | ( Ng853  &  (~ n2867) ) | ( (~ Ng1600)  &  (~ n2867) ) ;
 assign Ng30544 = ( (~ n2868) ) ;
 assign n2869 = ( (~ wire1594)  &  (~ Ng1597) ) | ( wire1594  &  (~ n2867) ) | ( (~ Ng1597)  &  (~ n2867) ) ;
 assign Ng30543 = ( (~ n2869) ) ;
 assign n2870 = ( (~ wire1612)  &  (~ Ng1594) ) | ( wire1612  &  (~ n2867) ) | ( (~ Ng1594)  &  (~ n2867) ) ;
 assign Ng30542 = ( (~ n2870) ) ;
 assign n2872 = ( (~ n1384)  &  n1469 ) | ( n1384  &  n3999 ) | ( n1469  &  n3999 ) ;
 assign n2873 = ( (~ Ng853)  &  (~ Ng1591) ) | ( Ng853  &  (~ n2872) ) | ( (~ Ng1591)  &  (~ n2872) ) ;
 assign Ng30541 = ( (~ n2873) ) ;
 assign n2874 = ( (~ wire1594)  &  (~ Ng1588) ) | ( wire1594  &  (~ n2872) ) | ( (~ Ng1588)  &  (~ n2872) ) ;
 assign Ng30540 = ( (~ n2874) ) ;
 assign n2875 = ( (~ wire1612)  &  (~ Ng1585) ) | ( wire1612  &  (~ n2872) ) | ( (~ Ng1585)  &  (~ n2872) ) ;
 assign Ng30539 = ( (~ n2875) ) ;
 assign n2877 = ( (~ n1384)  &  n1470 ) | ( n1384  &  n2711 ) | ( n1470  &  n2711 ) ;
 assign n2878 = ( (~ Ng853)  &  (~ Ng1573) ) | ( Ng853  &  (~ n2877) ) | ( (~ Ng1573)  &  (~ n2877) ) ;
 assign Ng30538 = ( (~ n2878) ) ;
 assign n2879 = ( (~ wire1594)  &  (~ Ng1570) ) | ( wire1594  &  (~ n2877) ) | ( (~ Ng1570)  &  (~ n2877) ) ;
 assign Ng30537 = ( (~ n2879) ) ;
 assign n2880 = ( (~ wire1612)  &  (~ Ng1567) ) | ( wire1612  &  (~ n2877) ) | ( (~ Ng1567)  &  (~ n2877) ) ;
 assign Ng30536 = ( (~ n2880) ) ;
 assign n2882 = ( (~ n1417)  &  n1475 ) | ( n1417  &  n4001 ) | ( n1475  &  n4001 ) ;
 assign n2883 = ( (~ Ng853)  &  (~ Ng951) ) | ( Ng853  &  (~ n2882) ) | ( (~ Ng951)  &  (~ n2882) ) ;
 assign Ng30535 = ( (~ n2883) ) ;
 assign n2884 = ( (~ wire1594)  &  (~ Ng948) ) | ( wire1594  &  (~ n2882) ) | ( (~ Ng948)  &  (~ n2882) ) ;
 assign Ng30534 = ( (~ n2884) ) ;
 assign n2885 = ( (~ wire1612)  &  (~ Ng945) ) | ( wire1612  &  (~ n2882) ) | ( (~ Ng945)  &  (~ n2882) ) ;
 assign Ng30533 = ( (~ n2885) ) ;
 assign n2886 = ( Ng853  &  n2124 ) | ( (~ Ng853)  &  (~ Ng942) ) | ( n2124  &  (~ Ng942) ) ;
 assign Ng30532 = ( (~ n2886) ) ;
 assign n2887 = ( wire1594  &  n2124 ) | ( (~ wire1594)  &  (~ Ng939) ) | ( n2124  &  (~ Ng939) ) ;
 assign Ng30531 = ( (~ n2887) ) ;
 assign n2888 = ( wire1612  &  n2124 ) | ( (~ wire1612)  &  (~ Ng936) ) | ( n2124  &  (~ Ng936) ) ;
 assign Ng30530 = ( (~ n2888) ) ;
 assign n2890 = ( (~ n1417)  &  n1476 ) | ( n1417  &  n4002 ) | ( n1476  &  n4002 ) ;
 assign n2891 = ( (~ Ng853)  &  (~ Ng906) ) | ( Ng853  &  (~ n2890) ) | ( (~ Ng906)  &  (~ n2890) ) ;
 assign Ng30529 = ( (~ n2891) ) ;
 assign n2892 = ( (~ wire1594)  &  (~ Ng903) ) | ( wire1594  &  (~ n2890) ) | ( (~ Ng903)  &  (~ n2890) ) ;
 assign Ng30528 = ( (~ n2892) ) ;
 assign n2893 = ( (~ wire1612)  &  (~ Ng900) ) | ( wire1612  &  (~ n2890) ) | ( (~ Ng900)  &  (~ n2890) ) ;
 assign Ng30527 = ( (~ n2893) ) ;
 assign n2895 = ( (~ n1417)  &  n1477 ) | ( n1417  &  n4003 ) | ( n1477  &  n4003 ) ;
 assign n2896 = ( (~ Ng853)  &  (~ Ng897) ) | ( Ng853  &  (~ n2895) ) | ( (~ Ng897)  &  (~ n2895) ) ;
 assign Ng30526 = ( (~ n2896) ) ;
 assign n2897 = ( (~ wire1594)  &  (~ Ng894) ) | ( wire1594  &  (~ n2895) ) | ( (~ Ng894)  &  (~ n2895) ) ;
 assign Ng30525 = ( (~ n2897) ) ;
 assign n2898 = ( (~ wire1612)  &  (~ Ng891) ) | ( wire1612  &  (~ n2895) ) | ( (~ Ng891)  &  (~ n2895) ) ;
 assign Ng30524 = ( (~ n2898) ) ;
 assign n2900 = ( (~ n1417)  &  n1478 ) | ( n1417  &  n2712 ) | ( n1478  &  n2712 ) ;
 assign n2901 = ( (~ Ng853)  &  (~ Ng879) ) | ( Ng853  &  (~ n2900) ) | ( (~ Ng879)  &  (~ n2900) ) ;
 assign Ng30523 = ( (~ n2901) ) ;
 assign n2902 = ( (~ wire1594)  &  (~ Ng876) ) | ( wire1594  &  (~ n2900) ) | ( (~ Ng876)  &  (~ n2900) ) ;
 assign Ng30522 = ( (~ n2902) ) ;
 assign n2903 = ( (~ wire1612)  &  (~ Ng873) ) | ( wire1612  &  (~ n2900) ) | ( (~ Ng873)  &  (~ n2900) ) ;
 assign Ng30521 = ( (~ n2903) ) ;
 assign n2905 = ( (~ n1450)  &  n1483 ) | ( n1450  &  n4005 ) | ( n1483  &  n4005 ) ;
 assign n2906 = ( (~ Ng853)  &  (~ Ng264) ) | ( Ng853  &  (~ n2905) ) | ( (~ Ng264)  &  (~ n2905) ) ;
 assign Ng30520 = ( (~ n2906) ) ;
 assign n2907 = ( (~ wire1594)  &  (~ Ng261) ) | ( wire1594  &  (~ n2905) ) | ( (~ Ng261)  &  (~ n2905) ) ;
 assign Ng30519 = ( (~ n2907) ) ;
 assign n2908 = ( (~ wire1612)  &  (~ Ng258) ) | ( wire1612  &  (~ n2905) ) | ( (~ Ng258)  &  (~ n2905) ) ;
 assign Ng30518 = ( (~ n2908) ) ;
 assign n2909 = ( Ng853  &  n2126 ) | ( (~ Ng853)  &  (~ Ng255) ) | ( n2126  &  (~ Ng255) ) ;
 assign Ng30517 = ( (~ n2909) ) ;
 assign n2910 = ( wire1594  &  n2126 ) | ( (~ wire1594)  &  (~ Ng252) ) | ( n2126  &  (~ Ng252) ) ;
 assign Ng30516 = ( (~ n2910) ) ;
 assign n2911 = ( wire1612  &  n2126 ) | ( (~ wire1612)  &  (~ Ng249) ) | ( n2126  &  (~ Ng249) ) ;
 assign Ng30515 = ( (~ n2911) ) ;
 assign n2913 = ( (~ n1450)  &  n1484 ) | ( n1450  &  n4006 ) | ( n1484  &  n4006 ) ;
 assign n2914 = ( (~ Ng853)  &  (~ Ng219) ) | ( Ng853  &  (~ n2913) ) | ( (~ Ng219)  &  (~ n2913) ) ;
 assign Ng30514 = ( (~ n2914) ) ;
 assign n2915 = ( (~ wire1594)  &  (~ Ng216) ) | ( wire1594  &  (~ n2913) ) | ( (~ Ng216)  &  (~ n2913) ) ;
 assign Ng30513 = ( (~ n2915) ) ;
 assign n2916 = ( (~ wire1612)  &  (~ Ng213) ) | ( wire1612  &  (~ n2913) ) | ( (~ Ng213)  &  (~ n2913) ) ;
 assign Ng30512 = ( (~ n2916) ) ;
 assign n2918 = ( (~ n1450)  &  n1485 ) | ( n1450  &  n4007 ) | ( n1485  &  n4007 ) ;
 assign n2919 = ( (~ Ng853)  &  (~ Ng210) ) | ( Ng853  &  (~ n2918) ) | ( (~ Ng210)  &  (~ n2918) ) ;
 assign Ng30511 = ( (~ n2919) ) ;
 assign n2920 = ( (~ wire1594)  &  (~ Ng207) ) | ( wire1594  &  (~ n2918) ) | ( (~ Ng207)  &  (~ n2918) ) ;
 assign Ng30510 = ( (~ n2920) ) ;
 assign n2921 = ( (~ wire1612)  &  (~ Ng204) ) | ( wire1612  &  (~ n2918) ) | ( (~ Ng204)  &  (~ n2918) ) ;
 assign Ng30509 = ( (~ n2921) ) ;
 assign n2923 = ( (~ n1450)  &  n1486 ) | ( n1450  &  n2713 ) | ( n1486  &  n2713 ) ;
 assign n2924 = ( (~ Ng853)  &  (~ Ng192) ) | ( Ng853  &  (~ n2923) ) | ( (~ Ng192)  &  (~ n2923) ) ;
 assign Ng30508 = ( (~ n2924) ) ;
 assign n2925 = ( (~ wire1594)  &  (~ Ng189) ) | ( wire1594  &  (~ n2923) ) | ( (~ Ng189)  &  (~ n2923) ) ;
 assign Ng30507 = ( (~ n2925) ) ;
 assign n2926 = ( (~ wire1612)  &  (~ Ng186) ) | ( wire1612  &  (~ n2923) ) | ( (~ Ng186)  &  (~ n2923) ) ;
 assign Ng30506 = ( (~ n2926) ) ;
 assign Ng29440 = ( n4013  &  (~ Ng1886) ) | ( n4013  &  Ng1887 ) | ( Ng1886  &  Ng1887 ) ;
 assign n2928 = ( n4016  &  (~ Ng2580) ) | ( n4016  &  (~ Ng2581) ) | ( Ng2580  &  (~ Ng2581) ) ;
 assign Ng30320 = ( (~ n2928) ) ;
 assign n2929 = ( wire1594  &  n4020 ) | ( (~ Ng305)  &  n4020 ) | ( (~ Ng299)  &  n4020 ) ;
 assign Ng23148 = ( (~ n2929) ) ;
 assign n2930 = ( n4022  &  Ng986 ) | ( n4022  &  Ng985 ) | ( (~ Ng986)  &  Ng985 ) ;
 assign Ng27200 = ( (~ n2930) ) ;
 assign n2931 = ( n4025  &  Ng1680 ) | ( n4025  &  Ng1679 ) | ( (~ Ng1680)  &  Ng1679 ) ;
 assign Ng29428 = ( (~ n2931) ) ;
 assign n2932 = ( n4028  &  Ng2374 ) | ( n4028  &  Ng2373 ) | ( (~ Ng2374)  &  Ng2373 ) ;
 assign Ng30314 = ( (~ n2932) ) ;
 assign n2933 = ( (~ Ng1315)  &  (~ Ng3105) ) | ( Ng1315  &  n2729 ) | ( (~ Ng3105)  &  n2729 ) ;
 assign Ng30122 = ( (~ n2933) ) ;
 assign n2934 = ( (~ wire1603)  &  (~ Ng3104) ) | ( wire1603  &  n2729 ) | ( (~ Ng3104)  &  n2729 ) ;
 assign Ng30121 = ( (~ n2934) ) ;
 assign n2935 = ( (~ wire1605)  &  (~ Ng3103) ) | ( wire1605  &  n2729 ) | ( (~ Ng3103)  &  n2729 ) ;
 assign Ng30120 = ( (~ n2935) ) ;
 assign n2936 = ( n515  &  (~ n557) ) | ( (~ n515)  &  (~ n1022) ) | ( (~ n557)  &  (~ n1022) ) ;
 assign n2937 = ( n256  &  (~ n654) ) | ( (~ n256)  &  n3739 ) | ( (~ n654)  &  n3739 ) ;
 assign n2938 = ( n282  &  (~ n654) ) | ( (~ n282)  &  n3739 ) | ( (~ n654)  &  n3739 ) ;
 assign n2939 = ( n358  &  (~ n654) ) | ( (~ n358)  &  n3739 ) | ( (~ n654)  &  n3739 ) ;
 assign n2940 = ( n317  &  (~ n557) ) | ( (~ n317)  &  (~ n1022) ) | ( (~ n557)  &  (~ n1022) ) ;
 assign n2941 = ( (~ Ng853)  &  (~ Ng2389) ) | ( Ng853  &  n4037 ) | ( (~ Ng2389)  &  n4037 ) ;
 assign Ng29809 = ( (~ n2941) ) ;
 assign n2942 = ( (~ wire1594)  &  (~ Ng2388) ) | ( wire1594  &  n4037 ) | ( (~ Ng2388)  &  n4037 ) ;
 assign Ng29808 = ( (~ n2942) ) ;
 assign n2943 = ( (~ wire1612)  &  (~ Ng2387) ) | ( wire1612  &  n4037 ) | ( (~ Ng2387)  &  n4037 ) ;
 assign Ng29807 = ( (~ n2943) ) ;
 assign n2944 = ( (~ Ng853)  &  (~ Ng1695) ) | ( Ng853  &  n4041 ) | ( (~ Ng1695)  &  n4041 ) ;
 assign Ng29805 = ( (~ n2944) ) ;
 assign n2945 = ( (~ wire1594)  &  (~ Ng1694) ) | ( wire1594  &  n4041 ) | ( (~ Ng1694)  &  n4041 ) ;
 assign Ng29804 = ( (~ n2945) ) ;
 assign n2946 = ( (~ wire1612)  &  (~ Ng1693) ) | ( wire1612  &  n4041 ) | ( (~ Ng1693)  &  n4041 ) ;
 assign Ng29803 = ( (~ n2946) ) ;
 assign n2947 = ( (~ Ng853)  &  (~ Ng1001) ) | ( Ng853  &  n4045 ) | ( (~ Ng1001)  &  n4045 ) ;
 assign Ng29801 = ( (~ n2947) ) ;
 assign n2948 = ( (~ wire1594)  &  (~ Ng1000) ) | ( wire1594  &  n4045 ) | ( (~ Ng1000)  &  n4045 ) ;
 assign Ng29800 = ( (~ n2948) ) ;
 assign n2949 = ( (~ wire1612)  &  (~ Ng999) ) | ( wire1612  &  n4045 ) | ( (~ Ng999)  &  n4045 ) ;
 assign Ng29799 = ( (~ n2949) ) ;
 assign n2950 = ( (~ Ng853)  &  (~ Ng314) ) | ( Ng853  &  n4049 ) | ( (~ Ng314)  &  n4049 ) ;
 assign Ng29797 = ( (~ n2950) ) ;
 assign n2951 = ( (~ wire1594)  &  (~ Ng313) ) | ( wire1594  &  n4049 ) | ( (~ Ng313)  &  n4049 ) ;
 assign Ng29796 = ( (~ n2951) ) ;
 assign n2952 = ( (~ wire1612)  &  (~ Ng312) ) | ( wire1612  &  n4049 ) | ( (~ Ng312)  &  n4049 ) ;
 assign Ng29795 = ( (~ n2952) ) ;
 assign n2954 = ( (~ Ng3147)  &  (~ n1768) ) | ( Ng3147  &  n1974 ) | ( (~ n1768)  &  n1974 ) ;
 assign n2955 = ( n493  &  (~ n548) ) | ( (~ n493)  &  (~ n993) ) | ( (~ n548)  &  (~ n993) ) ;
 assign n2956 = ( n228  &  (~ n649) ) | ( (~ n228)  &  n3738 ) | ( (~ n649)  &  n3738 ) ;
 assign n2957 = ( n247  &  (~ n649) ) | ( (~ n247)  &  n3738 ) | ( (~ n649)  &  n3738 ) ;
 assign n2958 = ( n308  &  (~ n649) ) | ( (~ n308)  &  n3738 ) | ( (~ n649)  &  n3738 ) ;
 assign n2959 = ( n275  &  (~ n548) ) | ( (~ n275)  &  (~ n993) ) | ( (~ n548)  &  (~ n993) ) ;
 assign n2960 = ( (~ Ng853)  &  (~ Ng2498) ) | ( Ng853  &  n4059 ) | ( (~ Ng2498)  &  n4059 ) ;
 assign Ng29654 = ( (~ n2960) ) ;
 assign n2961 = ( (~ wire1594)  &  (~ Ng2495) ) | ( wire1594  &  n4059 ) | ( (~ Ng2495)  &  n4059 ) ;
 assign Ng29653 = ( (~ n2961) ) ;
 assign n2962 = ( (~ wire1612)  &  (~ Ng2492) ) | ( wire1612  &  n4059 ) | ( (~ Ng2492)  &  n4059 ) ;
 assign Ng29652 = ( (~ n2962) ) ;
 assign n2963 = ( (~ n1542)  &  (~ Ng2396) ) | ( (~ n1542)  &  n4062 ) | ( (~ Ng2396)  &  (~ n4062) ) ;
 assign Ng29651 = ( (~ n2963) ) ;
 assign n2964 = ( (~ Ng2398)  &  (~ n1542) ) | ( (~ n1542)  &  n4066 ) | ( (~ Ng2398)  &  (~ n4066) ) ;
 assign Ng29650 = ( (~ n2964) ) ;
 assign n2965 = ( (~ n1542)  &  (~ Ng2397) ) | ( (~ n1542)  &  n4069 ) | ( (~ Ng2397)  &  (~ n4069) ) ;
 assign Ng29649 = ( (~ n2965) ) ;
 assign n2966 = ( (~ Ng853)  &  (~ Ng1804) ) | ( Ng853  &  n4071 ) | ( (~ Ng1804)  &  n4071 ) ;
 assign Ng29647 = ( (~ n2966) ) ;
 assign n2967 = ( (~ wire1594)  &  (~ Ng1801) ) | ( wire1594  &  n4071 ) | ( (~ Ng1801)  &  n4071 ) ;
 assign Ng29646 = ( (~ n2967) ) ;
 assign n2968 = ( (~ wire1612)  &  (~ Ng1798) ) | ( wire1612  &  n4071 ) | ( (~ Ng1798)  &  n4071 ) ;
 assign Ng29645 = ( (~ n2968) ) ;
 assign n2969 = ( (~ n1552)  &  (~ Ng1702) ) | ( (~ n1552)  &  n4074 ) | ( (~ Ng1702)  &  (~ n4074) ) ;
 assign Ng29644 = ( (~ n2969) ) ;
 assign n2970 = ( (~ Ng1704)  &  (~ n1552) ) | ( (~ n1552)  &  n4078 ) | ( (~ Ng1704)  &  (~ n4078) ) ;
 assign Ng29643 = ( (~ n2970) ) ;
 assign n2971 = ( (~ n1552)  &  (~ Ng1703) ) | ( (~ n1552)  &  n4081 ) | ( (~ Ng1703)  &  (~ n4081) ) ;
 assign Ng29642 = ( (~ n2971) ) ;
 assign n2972 = ( (~ Ng853)  &  (~ Ng1110) ) | ( Ng853  &  n4083 ) | ( (~ Ng1110)  &  n4083 ) ;
 assign Ng29640 = ( (~ n2972) ) ;
 assign n2973 = ( (~ wire1594)  &  (~ Ng1107) ) | ( wire1594  &  n4083 ) | ( (~ Ng1107)  &  n4083 ) ;
 assign Ng29639 = ( (~ n2973) ) ;
 assign n2974 = ( (~ wire1612)  &  (~ Ng1104) ) | ( wire1612  &  n4083 ) | ( (~ Ng1104)  &  n4083 ) ;
 assign Ng29638 = ( (~ n2974) ) ;
 assign n2975 = ( (~ n1562)  &  (~ Ng1008) ) | ( (~ n1562)  &  n4086 ) | ( (~ Ng1008)  &  (~ n4086) ) ;
 assign Ng29637 = ( (~ n2975) ) ;
 assign n2976 = ( (~ Ng1010)  &  (~ n1562) ) | ( (~ n1562)  &  n4090 ) | ( (~ Ng1010)  &  (~ n4090) ) ;
 assign Ng29636 = ( (~ n2976) ) ;
 assign n2977 = ( (~ n1562)  &  (~ Ng1009) ) | ( (~ n1562)  &  n4093 ) | ( (~ Ng1009)  &  (~ n4093) ) ;
 assign Ng29635 = ( (~ n2977) ) ;
 assign n2978 = ( (~ Ng853)  &  (~ Ng423) ) | ( Ng853  &  n4095 ) | ( (~ Ng423)  &  n4095 ) ;
 assign Ng29633 = ( (~ n2978) ) ;
 assign n2979 = ( (~ wire1594)  &  (~ Ng420) ) | ( wire1594  &  n4095 ) | ( (~ Ng420)  &  n4095 ) ;
 assign Ng29632 = ( (~ n2979) ) ;
 assign n2980 = ( (~ wire1612)  &  (~ Ng417) ) | ( wire1612  &  n4095 ) | ( (~ Ng417)  &  n4095 ) ;
 assign Ng29631 = ( (~ n2980) ) ;
 assign n2981 = ( (~ n1572)  &  (~ Ng321) ) | ( (~ n1572)  &  n4098 ) | ( (~ Ng321)  &  (~ n4098) ) ;
 assign Ng29630 = ( (~ n2981) ) ;
 assign n2982 = ( (~ Ng323)  &  (~ n1572) ) | ( (~ n1572)  &  n4102 ) | ( (~ Ng323)  &  (~ n4102) ) ;
 assign Ng29629 = ( (~ n2982) ) ;
 assign n2983 = ( (~ n1572)  &  (~ Ng322) ) | ( (~ n1572)  &  n4105 ) | ( (~ Ng322)  &  (~ n4105) ) ;
 assign Ng29628 = ( (~ n2983) ) ;
 assign n2984 = ( (~ Ng853)  &  (~ Ng2489) ) | ( Ng853  &  n4107 ) | ( (~ Ng2489)  &  n4107 ) ;
 assign Ng29449 = ( (~ n2984) ) ;
 assign n2985 = ( (~ wire1594)  &  (~ Ng2486) ) | ( wire1594  &  n4107 ) | ( (~ Ng2486)  &  n4107 ) ;
 assign Ng29448 = ( (~ n2985) ) ;
 assign n2986 = ( (~ wire1612)  &  (~ Ng2483) ) | ( wire1612  &  n4107 ) | ( (~ Ng2483)  &  n4107 ) ;
 assign Ng29447 = ( (~ n2986) ) ;
 assign n2987 = ( (~ Ng853)  &  (~ Ng1795) ) | ( Ng853  &  n4109 ) | ( (~ Ng1795)  &  n4109 ) ;
 assign Ng29436 = ( (~ n2987) ) ;
 assign n2988 = ( (~ wire1594)  &  (~ Ng1792) ) | ( wire1594  &  n4109 ) | ( (~ Ng1792)  &  n4109 ) ;
 assign Ng29435 = ( (~ n2988) ) ;
 assign n2989 = ( (~ wire1612)  &  (~ Ng1789) ) | ( wire1612  &  n4109 ) | ( (~ Ng1789)  &  n4109 ) ;
 assign Ng29434 = ( (~ n2989) ) ;
 assign n2990 = ( (~ Ng853)  &  (~ Ng1101) ) | ( Ng853  &  n4111 ) | ( (~ Ng1101)  &  n4111 ) ;
 assign Ng29423 = ( (~ n2990) ) ;
 assign n2991 = ( (~ wire1594)  &  (~ Ng1098) ) | ( wire1594  &  n4111 ) | ( (~ Ng1098)  &  n4111 ) ;
 assign Ng29422 = ( (~ n2991) ) ;
 assign n2992 = ( (~ wire1612)  &  (~ Ng1095) ) | ( wire1612  &  n4111 ) | ( (~ Ng1095)  &  n4111 ) ;
 assign Ng29421 = ( (~ n2992) ) ;
 assign n2993 = ( (~ Ng853)  &  (~ Ng414) ) | ( Ng853  &  n4113 ) | ( (~ Ng414)  &  n4113 ) ;
 assign Ng29416 = ( (~ n2993) ) ;
 assign n2994 = ( (~ wire1594)  &  (~ Ng411) ) | ( wire1594  &  n4113 ) | ( (~ Ng411)  &  n4113 ) ;
 assign Ng29415 = ( (~ n2994) ) ;
 assign n2995 = ( (~ wire1612)  &  (~ Ng408) ) | ( wire1612  &  n4113 ) | ( (~ Ng408)  &  n4113 ) ;
 assign Ng29414 = ( (~ n2995) ) ;
 assign n2996 = ( (~ Ng1315)  &  (~ Ng3102) ) | ( Ng1315  &  n2728 ) | ( (~ Ng3102)  &  n2728 ) ;
 assign Ng29165 = ( (~ n2996) ) ;
 assign n2997 = ( (~ wire1603)  &  (~ Ng3101) ) | ( wire1603  &  n2728 ) | ( (~ Ng3101)  &  n2728 ) ;
 assign Ng29164 = ( (~ n2997) ) ;
 assign n2998 = ( (~ wire1605)  &  (~ Ng3100) ) | ( wire1605  &  n2728 ) | ( (~ Ng3100)  &  n2728 ) ;
 assign Ng29163 = ( (~ n2998) ) ;
 assign n3000 = ( n109  &  (~ n1653) ) | ( (~ n103)  &  n109  &  (~ n1647) ) ;
 assign n3003 = ( n693  &  (~ n1656) ) | ( (~ n1656)  &  n1659 ) | ( n693  &  (~ n1659) ) ;
 assign n3004 = ( (~ Ng1315)  &  (~ Ng2694) ) | ( Ng1315  &  n4116 ) | ( (~ Ng2694)  &  n4116 ) ;
 assign Ng29161 = ( (~ n3004) ) ;
 assign n3005 = ( (~ wire1603)  &  (~ Ng2691) ) | ( wire1603  &  n4116 ) | ( (~ Ng2691)  &  n4116 ) ;
 assign Ng29160 = ( (~ n3005) ) ;
 assign n3006 = ( (~ wire1605)  &  (~ Ng2688) ) | ( wire1605  &  n4116 ) | ( (~ Ng2688)  &  n4116 ) ;
 assign Ng29159 = ( (~ n3006) ) ;
 assign n3008 = ( n693 ) | ( n1659 ) ;
 assign n3007 = ( (~ n693)  &  n1656  &  n3008 ) | ( n1656  &  n2545  &  n3008 ) ;
 assign n3009 = ( (~ Ng1315)  &  (~ Ng2685) ) | ( Ng1315  &  n4120 ) | ( (~ Ng2685)  &  n4120 ) ;
 assign Ng29158 = ( (~ n3009) ) ;
 assign n3010 = ( (~ wire1603)  &  (~ Ng2682) ) | ( wire1603  &  n4120 ) | ( (~ Ng2682)  &  n4120 ) ;
 assign Ng29157 = ( (~ n3010) ) ;
 assign n3011 = ( (~ wire1605)  &  (~ Ng2679) ) | ( wire1605  &  n4120 ) | ( (~ Ng2679)  &  n4120 ) ;
 assign Ng29156 = ( (~ n3011) ) ;
 assign n3013 = ( n100  &  (~ n1688) ) | ( (~ n91)  &  n100  &  (~ n1682) ) ;
 assign n3016 = ( n689  &  (~ n1691) ) | ( (~ n1691)  &  n1694 ) | ( n689  &  (~ n1694) ) ;
 assign n3017 = ( (~ Ng1315)  &  (~ Ng2000) ) | ( Ng1315  &  n4122 ) | ( (~ Ng2000)  &  n4122 ) ;
 assign Ng29153 = ( (~ n3017) ) ;
 assign n3018 = ( (~ wire1603)  &  (~ Ng1997) ) | ( wire1603  &  n4122 ) | ( (~ Ng1997)  &  n4122 ) ;
 assign Ng29152 = ( (~ n3018) ) ;
 assign n3019 = ( (~ wire1605)  &  (~ Ng1994) ) | ( wire1605  &  n4122 ) | ( (~ Ng1994)  &  n4122 ) ;
 assign Ng29151 = ( (~ n3019) ) ;
 assign n3021 = ( n689 ) | ( n1694 ) ;
 assign n3020 = ( (~ n689)  &  n1691  &  n3021 ) | ( n1691  &  n2571  &  n3021 ) ;
 assign n3022 = ( (~ Ng1315)  &  (~ Ng1991) ) | ( Ng1315  &  n4125 ) | ( (~ Ng1991)  &  n4125 ) ;
 assign Ng29150 = ( (~ n3022) ) ;
 assign n3023 = ( (~ wire1603)  &  (~ Ng1988) ) | ( wire1603  &  n4125 ) | ( (~ Ng1988)  &  n4125 ) ;
 assign Ng29149 = ( (~ n3023) ) ;
 assign n3024 = ( (~ wire1605)  &  (~ Ng1985) ) | ( wire1605  &  n4125 ) | ( (~ Ng1985)  &  n4125 ) ;
 assign Ng29148 = ( (~ n3024) ) ;
 assign n3026 = ( n88  &  (~ n1723) ) | ( (~ n79)  &  n88  &  (~ n1717) ) ;
 assign n3029 = ( n685  &  (~ n1726) ) | ( (~ n1726)  &  n1729 ) | ( n685  &  (~ n1729) ) ;
 assign n3030 = ( (~ Ng1315)  &  (~ Ng1306) ) | ( Ng1315  &  n4127 ) | ( (~ Ng1306)  &  n4127 ) ;
 assign Ng29145 = ( (~ n3030) ) ;
 assign n3031 = ( (~ wire1603)  &  (~ Ng1303) ) | ( wire1603  &  n4127 ) | ( (~ Ng1303)  &  n4127 ) ;
 assign Ng29144 = ( (~ n3031) ) ;
 assign n3032 = ( (~ wire1605)  &  (~ Ng1300) ) | ( wire1605  &  n4127 ) | ( (~ Ng1300)  &  n4127 ) ;
 assign Ng29143 = ( (~ n3032) ) ;
 assign n3034 = ( n685 ) | ( n1729 ) ;
 assign n3033 = ( (~ n685)  &  n1726  &  n3034 ) | ( n1726  &  n2595  &  n3034 ) ;
 assign n3035 = ( (~ Ng1315)  &  (~ Ng1297) ) | ( Ng1315  &  n4130 ) | ( (~ Ng1297)  &  n4130 ) ;
 assign Ng29142 = ( (~ n3035) ) ;
 assign n3036 = ( (~ wire1603)  &  (~ Ng1294) ) | ( wire1603  &  n4130 ) | ( (~ Ng1294)  &  n4130 ) ;
 assign Ng29141 = ( (~ n3036) ) ;
 assign n3037 = ( (~ wire1605)  &  (~ Ng1291) ) | ( wire1605  &  n4130 ) | ( (~ Ng1291)  &  n4130 ) ;
 assign Ng29140 = ( (~ n3037) ) ;
 assign n3039 = ( n76  &  (~ n1758) ) | ( (~ n70)  &  n76  &  (~ n1752) ) ;
 assign n3042 = ( n681  &  (~ n1761) ) | ( (~ n1761)  &  n1764 ) | ( n681  &  (~ n1764) ) ;
 assign n3043 = ( (~ Ng1315)  &  (~ Ng620) ) | ( Ng1315  &  n4132 ) | ( (~ Ng620)  &  n4132 ) ;
 assign Ng29137 = ( (~ n3043) ) ;
 assign n3044 = ( (~ wire1603)  &  (~ Ng617) ) | ( wire1603  &  n4132 ) | ( (~ Ng617)  &  n4132 ) ;
 assign Ng29136 = ( (~ n3044) ) ;
 assign n3045 = ( (~ wire1605)  &  (~ Ng614) ) | ( wire1605  &  n4132 ) | ( (~ Ng614)  &  n4132 ) ;
 assign Ng29135 = ( (~ n3045) ) ;
 assign n3047 = ( n681 ) | ( n1764 ) ;
 assign n3046 = ( (~ n681)  &  n1761  &  n3047 ) | ( n1761  &  n2619  &  n3047 ) ;
 assign n3048 = ( (~ Ng1315)  &  (~ Ng611) ) | ( Ng1315  &  n4135 ) | ( (~ Ng611)  &  n4135 ) ;
 assign Ng29134 = ( (~ n3048) ) ;
 assign n3049 = ( (~ wire1603)  &  (~ Ng608) ) | ( wire1603  &  n4135 ) | ( (~ Ng608)  &  n4135 ) ;
 assign Ng29133 = ( (~ n3049) ) ;
 assign n3050 = ( (~ wire1605)  &  (~ Ng605) ) | ( wire1605  &  n4135 ) | ( (~ Ng605)  &  n4135 ) ;
 assign Ng29132 = ( (~ n3050) ) ;
 assign n3051 = ( (~ Ng2658)  &  n4140 ) | ( (~ Ng2658)  &  n4142 ) | ( (~ n4140)  &  n4142 ) ;
 assign Ng28308 = ( (~ n3051) ) ;
 assign n3052 = ( (~ Ng2660)  &  n4142 ) | ( (~ Ng2660)  &  n4144 ) | ( n4142  &  (~ n4144) ) ;
 assign Ng28307 = ( (~ n3052) ) ;
 assign n3053 = ( (~ Ng2659)  &  n4142 ) | ( (~ Ng2659)  &  n4147 ) | ( n4142  &  (~ n4147) ) ;
 assign Ng28306 = ( (~ n3053) ) ;
 assign n3055 = ( n611  &  n2534 ) | ( n611  &  n4150 ) | ( n2534  &  (~ n4150) ) ;
 assign n3056 = ( (~ n3055)  &  (~ Ng2655) ) | ( (~ Ng2655)  &  n4140 ) | ( (~ n3055)  &  (~ n4140) ) ;
 assign Ng28305 = ( (~ n3056) ) ;
 assign n3057 = ( (~ Ng2657)  &  (~ n3055) ) | ( (~ Ng2657)  &  n4144 ) | ( (~ n3055)  &  (~ n4144) ) ;
 assign Ng28304 = ( (~ n3057) ) ;
 assign n3058 = ( (~ n3055)  &  (~ Ng2656) ) | ( (~ Ng2656)  &  n4147 ) | ( (~ n3055)  &  (~ n4147) ) ;
 assign Ng28303 = ( (~ n3058) ) ;
 assign n3060 = ( n611  &  n623 ) | ( n611  &  n4150 ) | ( (~ n623)  &  n4150 ) ;
 assign n3061 = ( (~ n3060)  &  (~ Ng2652) ) | ( (~ Ng2652)  &  n4140 ) | ( (~ n3060)  &  (~ n4140) ) ;
 assign Ng28302 = ( (~ n3061) ) ;
 assign n3062 = ( (~ Ng2654)  &  (~ n3060) ) | ( (~ Ng2654)  &  n4144 ) | ( (~ n3060)  &  (~ n4144) ) ;
 assign Ng28301 = ( (~ n3062) ) ;
 assign n3063 = ( (~ n3060)  &  (~ Ng2653) ) | ( (~ Ng2653)  &  n4147 ) | ( (~ n3060)  &  (~ n4147) ) ;
 assign Ng28300 = ( (~ n3063) ) ;
 assign n3064 = ( (~ n1831)  &  (~ Ng2649) ) | ( (~ Ng2649)  &  n4140 ) | ( (~ n1831)  &  (~ n4140) ) ;
 assign Ng28299 = ( (~ n3064) ) ;
 assign n3065 = ( (~ Ng2651)  &  (~ n1831) ) | ( (~ Ng2651)  &  n4144 ) | ( (~ n1831)  &  (~ n4144) ) ;
 assign Ng28298 = ( (~ n3065) ) ;
 assign n3066 = ( (~ n1831)  &  (~ Ng2650) ) | ( (~ Ng2650)  &  n4147 ) | ( (~ n1831)  &  (~ n4147) ) ;
 assign Ng28297 = ( (~ n3066) ) ;
 assign n3067 = ( (~ Ng11589)  &  (~ n4163) ) | ( (~ Ng11589)  &  n4165 ) | ( n4163  &  n4165 ) ;
 assign Ng28296 = ( (~ n3067) ) ;
 assign n3068 = ( (~ Ng11588)  &  n4165 ) | ( n4165  &  n4167 ) | ( (~ Ng11588)  &  (~ n4167) ) ;
 assign Ng28295 = ( (~ n3068) ) ;
 assign n3069 = ( (~ Ng11587)  &  n4165 ) | ( n4165  &  n4170 ) | ( (~ Ng11587)  &  (~ n4170) ) ;
 assign Ng28294 = ( (~ n3069) ) ;
 assign n3071 = ( n486  &  (~ n4904) ) | ( (~ n2138)  &  (~ n4904) ) ;
 assign n3072 = ( (~ n3071)  &  (~ Ng11586) ) | ( (~ n3071)  &  n4163 ) | ( (~ Ng11586)  &  (~ n4163) ) ;
 assign Ng28293 = ( (~ n3072) ) ;
 assign n3073 = ( (~ Ng11585)  &  (~ n3071) ) | ( (~ n3071)  &  n4167 ) | ( (~ Ng11585)  &  (~ n4167) ) ;
 assign Ng28292 = ( (~ n3073) ) ;
 assign n3074 = ( (~ n3071)  &  (~ Ng11584) ) | ( (~ n3071)  &  n4170 ) | ( (~ Ng11584)  &  (~ n4170) ) ;
 assign Ng28291 = ( (~ n3074) ) ;
 assign n3076 = ( n486  &  n509 ) | ( n486  &  n2138 ) | ( (~ n509)  &  n2138 ) ;
 assign n3077 = ( (~ n3076)  &  (~ Ng11583) ) | ( (~ n3076)  &  n4163 ) | ( (~ Ng11583)  &  (~ n4163) ) ;
 assign Ng28290 = ( (~ n3077) ) ;
 assign n3078 = ( (~ Ng11582)  &  (~ n3076) ) | ( (~ n3076)  &  n4167 ) | ( (~ Ng11582)  &  (~ n4167) ) ;
 assign Ng28289 = ( (~ n3078) ) ;
 assign n3079 = ( (~ n3076)  &  (~ Ng11581) ) | ( (~ n3076)  &  n4170 ) | ( (~ Ng11581)  &  (~ n4170) ) ;
 assign Ng28288 = ( (~ n3079) ) ;
 assign n3080 = ( (~ n1835)  &  (~ Ng11580) ) | ( (~ n1835)  &  n4163 ) | ( (~ Ng11580)  &  (~ n4163) ) ;
 assign Ng28287 = ( (~ n3080) ) ;
 assign n3081 = ( (~ Ng11579)  &  (~ n1835) ) | ( (~ n1835)  &  n4167 ) | ( (~ Ng11579)  &  (~ n4167) ) ;
 assign Ng28286 = ( (~ n3081) ) ;
 assign n3082 = ( (~ n1835)  &  (~ Ng11578) ) | ( (~ n1835)  &  n4170 ) | ( (~ Ng11578)  &  (~ n4170) ) ;
 assign Ng28285 = ( (~ n3082) ) ;
 assign n3083 = ( (~ Ng1964)  &  n4187 ) | ( (~ Ng1964)  &  n4189 ) | ( (~ n4187)  &  n4189 ) ;
 assign Ng28282 = ( (~ n3083) ) ;
 assign n3084 = ( (~ Ng1966)  &  n4189 ) | ( (~ Ng1966)  &  n4191 ) | ( n4189  &  (~ n4191) ) ;
 assign Ng28281 = ( (~ n3084) ) ;
 assign n3085 = ( (~ Ng1965)  &  n4189 ) | ( (~ Ng1965)  &  n4194 ) | ( n4189  &  (~ n4194) ) ;
 assign Ng28280 = ( (~ n3085) ) ;
 assign n3087 = ( n597  &  n2560 ) | ( n597  &  n4197 ) | ( n2560  &  (~ n4197) ) ;
 assign n3088 = ( (~ n3087)  &  (~ Ng1961) ) | ( (~ Ng1961)  &  n4187 ) | ( (~ n3087)  &  (~ n4187) ) ;
 assign Ng28279 = ( (~ n3088) ) ;
 assign n3089 = ( (~ Ng1963)  &  (~ n3087) ) | ( (~ Ng1963)  &  n4191 ) | ( (~ n3087)  &  (~ n4191) ) ;
 assign Ng28278 = ( (~ n3089) ) ;
 assign n3090 = ( (~ n3087)  &  (~ Ng1962) ) | ( (~ Ng1962)  &  n4194 ) | ( (~ n3087)  &  (~ n4194) ) ;
 assign Ng28277 = ( (~ n3090) ) ;
 assign n3092 = ( n597  &  n609 ) | ( n597  &  n4197 ) | ( (~ n609)  &  n4197 ) ;
 assign n3093 = ( (~ n3092)  &  (~ Ng1958) ) | ( (~ Ng1958)  &  n4187 ) | ( (~ n3092)  &  (~ n4187) ) ;
 assign Ng28276 = ( (~ n3093) ) ;
 assign n3094 = ( (~ Ng1960)  &  (~ n3092) ) | ( (~ Ng1960)  &  n4191 ) | ( (~ n3092)  &  (~ n4191) ) ;
 assign Ng28275 = ( (~ n3094) ) ;
 assign n3095 = ( (~ n3092)  &  (~ Ng1959) ) | ( (~ Ng1959)  &  n4194 ) | ( (~ n3092)  &  (~ n4194) ) ;
 assign Ng28274 = ( (~ n3095) ) ;
 assign n3096 = ( (~ n1841)  &  (~ Ng1955) ) | ( (~ Ng1955)  &  n4187 ) | ( (~ n1841)  &  (~ n4187) ) ;
 assign Ng28273 = ( (~ n3096) ) ;
 assign n3097 = ( (~ Ng1957)  &  (~ n1841) ) | ( (~ Ng1957)  &  n4191 ) | ( (~ n1841)  &  (~ n4191) ) ;
 assign Ng28272 = ( (~ n3097) ) ;
 assign n3098 = ( (~ n1841)  &  (~ Ng1956) ) | ( (~ Ng1956)  &  n4194 ) | ( (~ n1841)  &  (~ n4194) ) ;
 assign Ng28271 = ( (~ n3098) ) ;
 assign n3099 = ( (~ Ng11562)  &  (~ n4210) ) | ( (~ Ng11562)  &  n4212 ) | ( n4210  &  n4212 ) ;
 assign Ng28270 = ( (~ n3099) ) ;
 assign n3100 = ( (~ Ng11561)  &  n4212 ) | ( n4212  &  n4214 ) | ( (~ Ng11561)  &  (~ n4214) ) ;
 assign Ng28269 = ( (~ n3100) ) ;
 assign n3101 = ( (~ Ng11560)  &  n4212 ) | ( n4212  &  n4217 ) | ( (~ Ng11560)  &  (~ n4217) ) ;
 assign Ng28268 = ( (~ n3101) ) ;
 assign n3103 = ( n441  &  (~ n4905) ) | ( (~ n2139)  &  (~ n4905) ) ;
 assign n3104 = ( (~ n3103)  &  (~ Ng11559) ) | ( (~ n3103)  &  n4210 ) | ( (~ Ng11559)  &  (~ n4210) ) ;
 assign Ng28267 = ( (~ n3104) ) ;
 assign n3105 = ( (~ Ng11558)  &  (~ n3103) ) | ( (~ n3103)  &  n4214 ) | ( (~ Ng11558)  &  (~ n4214) ) ;
 assign Ng28266 = ( (~ n3105) ) ;
 assign n3106 = ( (~ n3103)  &  (~ Ng11557) ) | ( (~ n3103)  &  n4217 ) | ( (~ Ng11557)  &  (~ n4217) ) ;
 assign Ng28265 = ( (~ n3106) ) ;
 assign n3108 = ( n441  &  n474 ) | ( n441  &  n2139 ) | ( (~ n474)  &  n2139 ) ;
 assign n3109 = ( (~ n3108)  &  (~ Ng11556) ) | ( (~ n3108)  &  n4210 ) | ( (~ Ng11556)  &  (~ n4210) ) ;
 assign Ng28264 = ( (~ n3109) ) ;
 assign n3110 = ( (~ Ng11555)  &  (~ n3108) ) | ( (~ n3108)  &  n4214 ) | ( (~ Ng11555)  &  (~ n4214) ) ;
 assign Ng28263 = ( (~ n3110) ) ;
 assign n3111 = ( (~ n3108)  &  (~ Ng11554) ) | ( (~ n3108)  &  n4217 ) | ( (~ Ng11554)  &  (~ n4217) ) ;
 assign Ng28262 = ( (~ n3111) ) ;
 assign n3112 = ( (~ n1844)  &  (~ Ng11553) ) | ( (~ n1844)  &  n4210 ) | ( (~ Ng11553)  &  (~ n4210) ) ;
 assign Ng28261 = ( (~ n3112) ) ;
 assign n3113 = ( (~ Ng11552)  &  (~ n1844) ) | ( (~ n1844)  &  n4214 ) | ( (~ Ng11552)  &  (~ n4214) ) ;
 assign Ng28260 = ( (~ n3113) ) ;
 assign n3114 = ( (~ n1844)  &  (~ Ng11551) ) | ( (~ n1844)  &  n4217 ) | ( (~ Ng11551)  &  (~ n4217) ) ;
 assign Ng28259 = ( (~ n3114) ) ;
 assign n3115 = ( (~ Ng1270)  &  n4234 ) | ( (~ Ng1270)  &  n4236 ) | ( (~ n4234)  &  n4236 ) ;
 assign Ng28256 = ( (~ n3115) ) ;
 assign n3116 = ( (~ Ng1272)  &  n4236 ) | ( (~ Ng1272)  &  n4238 ) | ( n4236  &  (~ n4238) ) ;
 assign Ng28255 = ( (~ n3116) ) ;
 assign n3117 = ( (~ Ng1271)  &  n4236 ) | ( (~ Ng1271)  &  n4241 ) | ( n4236  &  (~ n4241) ) ;
 assign Ng28254 = ( (~ n3117) ) ;
 assign n3119 = ( n583  &  n2584 ) | ( n583  &  n4244 ) | ( n2584  &  (~ n4244) ) ;
 assign n3120 = ( (~ n3119)  &  (~ Ng1267) ) | ( (~ Ng1267)  &  n4234 ) | ( (~ n3119)  &  (~ n4234) ) ;
 assign Ng28253 = ( (~ n3120) ) ;
 assign n3121 = ( (~ Ng1269)  &  (~ n3119) ) | ( (~ Ng1269)  &  n4238 ) | ( (~ n3119)  &  (~ n4238) ) ;
 assign Ng28252 = ( (~ n3121) ) ;
 assign n3122 = ( (~ n3119)  &  (~ Ng1268) ) | ( (~ Ng1268)  &  n4241 ) | ( (~ n3119)  &  (~ n4241) ) ;
 assign Ng28251 = ( (~ n3122) ) ;
 assign n3124 = ( n583  &  n595 ) | ( n583  &  n4244 ) | ( (~ n595)  &  n4244 ) ;
 assign n3125 = ( (~ n3124)  &  (~ Ng1264) ) | ( (~ Ng1264)  &  n4234 ) | ( (~ n3124)  &  (~ n4234) ) ;
 assign Ng28250 = ( (~ n3125) ) ;
 assign n3126 = ( (~ Ng1266)  &  (~ n3124) ) | ( (~ Ng1266)  &  n4238 ) | ( (~ n3124)  &  (~ n4238) ) ;
 assign Ng28249 = ( (~ n3126) ) ;
 assign n3127 = ( (~ n3124)  &  (~ Ng1265) ) | ( (~ Ng1265)  &  n4241 ) | ( (~ n3124)  &  (~ n4241) ) ;
 assign Ng28248 = ( (~ n3127) ) ;
 assign n3128 = ( (~ n1850)  &  (~ Ng1261) ) | ( (~ Ng1261)  &  n4234 ) | ( (~ n1850)  &  (~ n4234) ) ;
 assign Ng28247 = ( (~ n3128) ) ;
 assign n3129 = ( (~ Ng1263)  &  (~ n1850) ) | ( (~ Ng1263)  &  n4238 ) | ( (~ n1850)  &  (~ n4238) ) ;
 assign Ng28246 = ( (~ n3129) ) ;
 assign n3130 = ( (~ n1850)  &  (~ Ng1262) ) | ( (~ Ng1262)  &  n4241 ) | ( (~ n1850)  &  (~ n4241) ) ;
 assign Ng28245 = ( (~ n3130) ) ;
 assign n3131 = ( (~ Ng11535)  &  (~ n4257) ) | ( (~ Ng11535)  &  n4259 ) | ( n4257  &  n4259 ) ;
 assign Ng28244 = ( (~ n3131) ) ;
 assign n3132 = ( (~ Ng11534)  &  n4259 ) | ( n4259  &  n4261 ) | ( (~ Ng11534)  &  (~ n4261) ) ;
 assign Ng28243 = ( (~ n3132) ) ;
 assign n3133 = ( (~ Ng11533)  &  n4259 ) | ( n4259  &  n4264 ) | ( (~ Ng11533)  &  (~ n4264) ) ;
 assign Ng28242 = ( (~ n3133) ) ;
 assign n3135 = ( n391  &  (~ n4906) ) | ( (~ n2140)  &  (~ n4906) ) ;
 assign n3136 = ( (~ n3135)  &  (~ Ng11532) ) | ( (~ n3135)  &  n4257 ) | ( (~ Ng11532)  &  (~ n4257) ) ;
 assign Ng28241 = ( (~ n3136) ) ;
 assign n3137 = ( (~ Ng11531)  &  (~ n3135) ) | ( (~ n3135)  &  n4261 ) | ( (~ Ng11531)  &  (~ n4261) ) ;
 assign Ng28240 = ( (~ n3137) ) ;
 assign n3138 = ( (~ n3135)  &  (~ Ng11530) ) | ( (~ n3135)  &  n4264 ) | ( (~ Ng11530)  &  (~ n4264) ) ;
 assign Ng28239 = ( (~ n3138) ) ;
 assign n3140 = ( n391  &  n429 ) | ( n391  &  n2140 ) | ( (~ n429)  &  n2140 ) ;
 assign n3141 = ( (~ n3140)  &  (~ Ng11529) ) | ( (~ n3140)  &  n4257 ) | ( (~ Ng11529)  &  (~ n4257) ) ;
 assign Ng28238 = ( (~ n3141) ) ;
 assign n3142 = ( (~ Ng11528)  &  (~ n3140) ) | ( (~ n3140)  &  n4261 ) | ( (~ Ng11528)  &  (~ n4261) ) ;
 assign Ng28237 = ( (~ n3142) ) ;
 assign n3143 = ( (~ n3140)  &  (~ Ng11527) ) | ( (~ n3140)  &  n4264 ) | ( (~ Ng11527)  &  (~ n4264) ) ;
 assign Ng28236 = ( (~ n3143) ) ;
 assign n3144 = ( (~ n1853)  &  (~ Ng11526) ) | ( (~ n1853)  &  n4257 ) | ( (~ Ng11526)  &  (~ n4257) ) ;
 assign Ng28235 = ( (~ n3144) ) ;
 assign n3145 = ( (~ Ng11525)  &  (~ n1853) ) | ( (~ n1853)  &  n4261 ) | ( (~ Ng11525)  &  (~ n4261) ) ;
 assign Ng28234 = ( (~ n3145) ) ;
 assign n3146 = ( (~ n1853)  &  (~ Ng11524) ) | ( (~ n1853)  &  n4264 ) | ( (~ Ng11524)  &  (~ n4264) ) ;
 assign Ng28233 = ( (~ n3146) ) ;
 assign n3147 = ( (~ Ng584)  &  n4281 ) | ( (~ Ng584)  &  n4283 ) | ( (~ n4281)  &  n4283 ) ;
 assign Ng28230 = ( (~ n3147) ) ;
 assign n3148 = ( (~ Ng586)  &  n4283 ) | ( (~ Ng586)  &  n4285 ) | ( n4283  &  (~ n4285) ) ;
 assign Ng28229 = ( (~ n3148) ) ;
 assign n3149 = ( (~ Ng585)  &  n4283 ) | ( (~ Ng585)  &  n4288 ) | ( n4283  &  (~ n4288) ) ;
 assign Ng28228 = ( (~ n3149) ) ;
 assign n3151 = ( n574  &  n2608 ) | ( n574  &  n4291 ) | ( n2608  &  (~ n4291) ) ;
 assign n3152 = ( (~ n3151)  &  (~ Ng581) ) | ( (~ Ng581)  &  n4281 ) | ( (~ n3151)  &  (~ n4281) ) ;
 assign Ng28227 = ( (~ n3152) ) ;
 assign n3153 = ( (~ Ng583)  &  (~ n3151) ) | ( (~ Ng583)  &  n4285 ) | ( (~ n3151)  &  (~ n4285) ) ;
 assign Ng28226 = ( (~ n3153) ) ;
 assign n3154 = ( (~ n3151)  &  (~ Ng582) ) | ( (~ Ng582)  &  n4288 ) | ( (~ n3151)  &  (~ n4288) ) ;
 assign Ng28225 = ( (~ n3154) ) ;
 assign n3156 = ( n574  &  n581 ) | ( n574  &  n4291 ) | ( (~ n581)  &  n4291 ) ;
 assign n3157 = ( (~ n3156)  &  (~ Ng578) ) | ( (~ Ng578)  &  n4281 ) | ( (~ n3156)  &  (~ n4281) ) ;
 assign Ng28224 = ( (~ n3157) ) ;
 assign n3158 = ( (~ Ng580)  &  (~ n3156) ) | ( (~ Ng580)  &  n4285 ) | ( (~ n3156)  &  (~ n4285) ) ;
 assign Ng28223 = ( (~ n3158) ) ;
 assign n3159 = ( (~ n3156)  &  (~ Ng579) ) | ( (~ Ng579)  &  n4288 ) | ( (~ n3156)  &  (~ n4288) ) ;
 assign Ng28222 = ( (~ n3159) ) ;
 assign n3160 = ( (~ n1859)  &  (~ Ng575) ) | ( (~ Ng575)  &  n4281 ) | ( (~ n1859)  &  (~ n4281) ) ;
 assign Ng28221 = ( (~ n3160) ) ;
 assign n3161 = ( (~ Ng577)  &  (~ n1859) ) | ( (~ Ng577)  &  n4285 ) | ( (~ n1859)  &  (~ n4285) ) ;
 assign Ng28220 = ( (~ n3161) ) ;
 assign n3162 = ( (~ n1859)  &  (~ Ng576) ) | ( (~ Ng576)  &  n4288 ) | ( (~ n1859)  &  (~ n4288) ) ;
 assign Ng28219 = ( (~ n3162) ) ;
 assign n3163 = ( (~ Ng11508)  &  (~ n4304) ) | ( (~ Ng11508)  &  n4306 ) | ( n4304  &  n4306 ) ;
 assign Ng28218 = ( (~ n3163) ) ;
 assign n3164 = ( (~ Ng11507)  &  n4306 ) | ( n4306  &  n4308 ) | ( (~ Ng11507)  &  (~ n4308) ) ;
 assign Ng28217 = ( (~ n3164) ) ;
 assign n3165 = ( (~ Ng11506)  &  n4306 ) | ( n4306  &  n4311 ) | ( (~ Ng11506)  &  (~ n4311) ) ;
 assign Ng28216 = ( (~ n3165) ) ;
 assign n3167 = ( n341  &  (~ n4907) ) | ( (~ n2141)  &  (~ n4907) ) ;
 assign n3168 = ( (~ n3167)  &  (~ Ng11505) ) | ( (~ n3167)  &  n4304 ) | ( (~ Ng11505)  &  (~ n4304) ) ;
 assign Ng28215 = ( (~ n3168) ) ;
 assign n3169 = ( (~ Ng11504)  &  (~ n3167) ) | ( (~ n3167)  &  n4308 ) | ( (~ Ng11504)  &  (~ n4308) ) ;
 assign Ng28214 = ( (~ n3169) ) ;
 assign n3170 = ( (~ n3167)  &  (~ Ng11503) ) | ( (~ n3167)  &  n4311 ) | ( (~ Ng11503)  &  (~ n4311) ) ;
 assign Ng28213 = ( (~ n3170) ) ;
 assign n3172 = ( n341  &  n379 ) | ( n341  &  n2141 ) | ( (~ n379)  &  n2141 ) ;
 assign n3173 = ( (~ n3172)  &  (~ Ng11502) ) | ( (~ n3172)  &  n4304 ) | ( (~ Ng11502)  &  (~ n4304) ) ;
 assign Ng28212 = ( (~ n3173) ) ;
 assign n3174 = ( (~ Ng11501)  &  (~ n3172) ) | ( (~ n3172)  &  n4308 ) | ( (~ Ng11501)  &  (~ n4308) ) ;
 assign Ng28211 = ( (~ n3174) ) ;
 assign n3175 = ( (~ n3172)  &  (~ Ng11500) ) | ( (~ n3172)  &  n4311 ) | ( (~ Ng11500)  &  (~ n4311) ) ;
 assign Ng28210 = ( (~ n3175) ) ;
 assign n3176 = ( (~ n1862)  &  (~ Ng11499) ) | ( (~ n1862)  &  n4304 ) | ( (~ Ng11499)  &  (~ n4304) ) ;
 assign Ng28209 = ( (~ n3176) ) ;
 assign n3177 = ( (~ Ng11498)  &  (~ n1862) ) | ( (~ n1862)  &  n4308 ) | ( (~ Ng11498)  &  (~ n4308) ) ;
 assign Ng28208 = ( (~ n3177) ) ;
 assign n3178 = ( (~ n1862)  &  (~ Ng11497) ) | ( (~ n1862)  &  n4311 ) | ( (~ Ng11497)  &  (~ n4311) ) ;
 assign Ng28207 = ( (~ n3178) ) ;
 assign n3179 = ( (~ Ng853)  &  (~ Ng2519) ) | ( Ng853  &  n4328 ) | ( (~ Ng2519)  &  n4328 ) ;
 assign Ng27713 = ( (~ n3179) ) ;
 assign n3180 = ( (~ wire1594)  &  (~ Ng2516) ) | ( wire1594  &  n4328 ) | ( (~ Ng2516)  &  n4328 ) ;
 assign Ng27712 = ( (~ n3180) ) ;
 assign n3181 = ( (~ wire1612)  &  (~ Ng2513) ) | ( wire1612  &  n4328 ) | ( (~ Ng2513)  &  n4328 ) ;
 assign Ng27711 = ( (~ n3181) ) ;
 assign n3182 = ( (~ Ng853)  &  (~ Ng2510) ) | ( Ng853  &  n4329 ) | ( (~ Ng2510)  &  n4329 ) ;
 assign Ng27710 = ( (~ n3182) ) ;
 assign n3183 = ( (~ wire1594)  &  (~ Ng2507) ) | ( wire1594  &  n4329 ) | ( (~ Ng2507)  &  n4329 ) ;
 assign Ng27709 = ( (~ n3183) ) ;
 assign n3184 = ( (~ wire1612)  &  (~ Ng2504) ) | ( wire1612  &  n4329 ) | ( (~ Ng2504)  &  n4329 ) ;
 assign Ng27708 = ( (~ n3184) ) ;
 assign n3185 = ( (~ Ng853)  &  (~ Ng1825) ) | ( Ng853  &  n4330 ) | ( (~ Ng1825)  &  n4330 ) ;
 assign Ng27705 = ( (~ n3185) ) ;
 assign n3186 = ( (~ wire1594)  &  (~ Ng1822) ) | ( wire1594  &  n4330 ) | ( (~ Ng1822)  &  n4330 ) ;
 assign Ng27704 = ( (~ n3186) ) ;
 assign n3187 = ( (~ wire1612)  &  (~ Ng1819) ) | ( wire1612  &  n4330 ) | ( (~ Ng1819)  &  n4330 ) ;
 assign Ng27703 = ( (~ n3187) ) ;
 assign n3188 = ( (~ Ng853)  &  (~ Ng1816) ) | ( Ng853  &  n4331 ) | ( (~ Ng1816)  &  n4331 ) ;
 assign Ng27702 = ( (~ n3188) ) ;
 assign n3189 = ( (~ wire1594)  &  (~ Ng1813) ) | ( wire1594  &  n4331 ) | ( (~ Ng1813)  &  n4331 ) ;
 assign Ng27701 = ( (~ n3189) ) ;
 assign n3190 = ( (~ wire1612)  &  (~ Ng1810) ) | ( wire1612  &  n4331 ) | ( (~ Ng1810)  &  n4331 ) ;
 assign Ng27700 = ( (~ n3190) ) ;
 assign n3191 = ( (~ Ng853)  &  (~ Ng1131) ) | ( Ng853  &  n4332 ) | ( (~ Ng1131)  &  n4332 ) ;
 assign Ng27697 = ( (~ n3191) ) ;
 assign n3192 = ( (~ wire1594)  &  (~ Ng1128) ) | ( wire1594  &  n4332 ) | ( (~ Ng1128)  &  n4332 ) ;
 assign Ng27696 = ( (~ n3192) ) ;
 assign n3193 = ( (~ wire1612)  &  (~ Ng1125) ) | ( wire1612  &  n4332 ) | ( (~ Ng1125)  &  n4332 ) ;
 assign Ng27695 = ( (~ n3193) ) ;
 assign n3194 = ( (~ Ng853)  &  (~ Ng1122) ) | ( Ng853  &  n4333 ) | ( (~ Ng1122)  &  n4333 ) ;
 assign Ng27694 = ( (~ n3194) ) ;
 assign n3195 = ( (~ wire1594)  &  (~ Ng1119) ) | ( wire1594  &  n4333 ) | ( (~ Ng1119)  &  n4333 ) ;
 assign Ng27693 = ( (~ n3195) ) ;
 assign n3196 = ( (~ wire1612)  &  (~ Ng1116) ) | ( wire1612  &  n4333 ) | ( (~ Ng1116)  &  n4333 ) ;
 assign Ng27692 = ( (~ n3196) ) ;
 assign n3197 = ( (~ Ng853)  &  (~ Ng444) ) | ( Ng853  &  n4334 ) | ( (~ Ng444)  &  n4334 ) ;
 assign Ng27689 = ( (~ n3197) ) ;
 assign n3198 = ( (~ wire1594)  &  (~ Ng441) ) | ( wire1594  &  n4334 ) | ( (~ Ng441)  &  n4334 ) ;
 assign Ng27688 = ( (~ n3198) ) ;
 assign n3199 = ( (~ wire1612)  &  (~ Ng438) ) | ( wire1612  &  n4334 ) | ( (~ Ng438)  &  n4334 ) ;
 assign Ng27687 = ( (~ n3199) ) ;
 assign n3200 = ( (~ Ng853)  &  (~ Ng435) ) | ( Ng853  &  n4335 ) | ( (~ Ng435)  &  n4335 ) ;
 assign Ng27686 = ( (~ n3200) ) ;
 assign n3201 = ( (~ wire1594)  &  (~ Ng432) ) | ( wire1594  &  n4335 ) | ( (~ Ng432)  &  n4335 ) ;
 assign Ng27685 = ( (~ n3201) ) ;
 assign n3202 = ( (~ wire1612)  &  (~ Ng429) ) | ( wire1612  &  n4335 ) | ( (~ Ng429)  &  n4335 ) ;
 assign Ng27684 = ( (~ n3202) ) ;
 assign n3203 = ( (~ Ng1315)  &  (~ Ng2571) ) | ( Ng1315  &  n4336 ) | ( (~ Ng2571)  &  n4336 ) ;
 assign Ng27235 = ( (~ n3203) ) ;
 assign n3204 = ( (~ wire1603)  &  (~ Ng2568) ) | ( wire1603  &  n4336 ) | ( (~ Ng2568)  &  n4336 ) ;
 assign Ng27234 = ( (~ n3204) ) ;
 assign n3205 = ( (~ wire1605)  &  (~ Ng2565) ) | ( wire1605  &  n4336 ) | ( (~ Ng2565)  &  n4336 ) ;
 assign Ng27233 = ( (~ n3205) ) ;
 assign n3206 = ( (~ Ng2477)  &  n4337 ) | ( (~ Ng2477)  &  n4339 ) | ( (~ n4337)  &  n4339 ) ;
 assign Ng27232 = ( (~ n3206) ) ;
 assign n3207 = ( (~ Ng2479)  &  n4339 ) | ( (~ Ng2479)  &  n4341 ) | ( n4339  &  (~ n4341) ) ;
 assign Ng27231 = ( (~ n3207) ) ;
 assign n3208 = ( (~ Ng2478)  &  n4339 ) | ( (~ Ng2478)  &  n4344 ) | ( n4339  &  (~ n4344) ) ;
 assign Ng27230 = ( (~ n3208) ) ;
 assign n3209 = ( (~ Ng1315)  &  (~ Ng1877) ) | ( Ng1315  &  n4347 ) | ( (~ Ng1877)  &  n4347 ) ;
 assign Ng27226 = ( (~ n3209) ) ;
 assign n3210 = ( (~ wire1603)  &  (~ Ng1874) ) | ( wire1603  &  n4347 ) | ( (~ Ng1874)  &  n4347 ) ;
 assign Ng27225 = ( (~ n3210) ) ;
 assign n3211 = ( (~ wire1605)  &  (~ Ng1871) ) | ( wire1605  &  n4347 ) | ( (~ Ng1871)  &  n4347 ) ;
 assign Ng27224 = ( (~ n3211) ) ;
 assign n3212 = ( (~ Ng1783)  &  n4337 ) | ( (~ Ng1783)  &  n4349 ) | ( (~ n4337)  &  n4349 ) ;
 assign Ng27223 = ( (~ n3212) ) ;
 assign n3213 = ( (~ Ng1785)  &  n4341 ) | ( (~ Ng1785)  &  n4349 ) | ( (~ n4341)  &  n4349 ) ;
 assign Ng27222 = ( (~ n3213) ) ;
 assign n3214 = ( (~ Ng1784)  &  n4344 ) | ( (~ Ng1784)  &  n4349 ) | ( (~ n4344)  &  n4349 ) ;
 assign Ng27221 = ( (~ n3214) ) ;
 assign n3215 = ( (~ Ng1315)  &  (~ Ng1183) ) | ( Ng1315  &  n4352 ) | ( (~ Ng1183)  &  n4352 ) ;
 assign Ng27211 = ( (~ n3215) ) ;
 assign n3216 = ( (~ wire1603)  &  (~ Ng1180) ) | ( wire1603  &  n4352 ) | ( (~ Ng1180)  &  n4352 ) ;
 assign Ng27210 = ( (~ n3216) ) ;
 assign n3217 = ( (~ wire1605)  &  (~ Ng1177) ) | ( wire1605  &  n4352 ) | ( (~ Ng1177)  &  n4352 ) ;
 assign Ng27209 = ( (~ n3217) ) ;
 assign n3218 = ( (~ Ng1089)  &  n4337 ) | ( (~ Ng1089)  &  n4354 ) | ( (~ n4337)  &  n4354 ) ;
 assign Ng27208 = ( (~ n3218) ) ;
 assign n3219 = ( (~ Ng1091)  &  n4341 ) | ( (~ Ng1091)  &  n4354 ) | ( (~ n4341)  &  n4354 ) ;
 assign Ng27207 = ( (~ n3219) ) ;
 assign n3220 = ( (~ Ng1090)  &  n4344 ) | ( (~ Ng1090)  &  n4354 ) | ( (~ n4344)  &  n4354 ) ;
 assign Ng27206 = ( (~ n3220) ) ;
 assign n3221 = ( (~ Ng1315)  &  (~ Ng496) ) | ( Ng1315  &  n4357 ) | ( (~ Ng496)  &  n4357 ) ;
 assign Ng27196 = ( (~ n3221) ) ;
 assign n3222 = ( (~ wire1603)  &  (~ Ng493) ) | ( wire1603  &  n4357 ) | ( (~ Ng493)  &  n4357 ) ;
 assign Ng27195 = ( (~ n3222) ) ;
 assign n3223 = ( (~ wire1605)  &  (~ Ng490) ) | ( wire1605  &  n4357 ) | ( (~ Ng490)  &  n4357 ) ;
 assign Ng27194 = ( (~ n3223) ) ;
 assign n3224 = ( (~ Ng402)  &  n4337 ) | ( (~ Ng402)  &  n4359 ) | ( (~ n4337)  &  n4359 ) ;
 assign Ng27193 = ( (~ n3224) ) ;
 assign n3225 = ( (~ Ng404)  &  n4341 ) | ( (~ Ng404)  &  n4359 ) | ( (~ n4341)  &  n4359 ) ;
 assign Ng27192 = ( (~ n3225) ) ;
 assign n3226 = ( (~ Ng403)  &  n4344 ) | ( (~ Ng403)  &  n4359 ) | ( (~ n4344)  &  n4359 ) ;
 assign Ng27191 = ( (~ n3226) ) ;
 assign n3227 = ( (~ Ng1315)  &  (~ Ng3099) ) | ( Ng1315  &  n2727 ) | ( (~ Ng3099)  &  n2727 ) ;
 assign Ng26753 = ( (~ n3227) ) ;
 assign n3228 = ( (~ wire1603)  &  (~ Ng3098) ) | ( wire1603  &  n2727 ) | ( (~ Ng3098)  &  n2727 ) ;
 assign Ng26752 = ( (~ n3228) ) ;
 assign n3229 = ( (~ wire1605)  &  (~ Ng3097) ) | ( wire1605  &  n2727 ) | ( (~ Ng3097)  &  n2727 ) ;
 assign Ng26751 = ( (~ n3229) ) ;
 assign n3230 = ( Pg3234  &  n1905 ) | ( Pg3234  &  n4362 ) | ( (~ n1905)  &  n4362 ) ;
 assign Ng26748 = ( (~ n3230) ) ;
 assign n3231 = ( (~ n768)  &  n770 ) | ( (~ n768)  &  (~ Ng2808) ) | ( (~ n770)  &  (~ Ng2808) ) ;
 assign Ng26745 = ( (~ n3231) ) ;
 assign n3232 = ( n767  &  (~ n768) ) | ( (~ n767)  &  (~ Ng2810) ) | ( (~ n768)  &  (~ Ng2810) ) ;
 assign Ng26744 = ( (~ n3232) ) ;
 assign n3233 = ( n761  &  (~ n768) ) | ( (~ n761)  &  (~ Ng2809) ) | ( (~ n768)  &  (~ Ng2809) ) ;
 assign Ng26743 = ( (~ n3233) ) ;
 assign n3234 = ( n1789  &  (~ Ng2253) ) | ( (~ Ng2253)  &  n4370 ) | ( n1789  &  (~ n4370) ) ;
 assign Ng26741 = ( (~ n3234) ) ;
 assign n3235 = ( n1789  &  (~ n4373) ) | ( n1789  &  (~ Ng2255) ) | ( n4373  &  (~ Ng2255) ) ;
 assign Ng26740 = ( (~ n3235) ) ;
 assign n3236 = ( n1789  &  (~ Ng2254) ) | ( (~ Ng2254)  &  n4375 ) | ( n1789  &  (~ n4375) ) ;
 assign Ng26739 = ( (~ n3236) ) ;
 assign n3237 = ( Ng2165  &  (~ Ng2250) ) | ( (~ Ng2250)  &  n4370 ) | ( Ng2165  &  (~ n4370) ) ;
 assign Ng26738 = ( (~ n3237) ) ;
 assign n3238 = ( (~ Ng2252)  &  Ng2165 ) | ( (~ Ng2252)  &  n4373 ) | ( Ng2165  &  (~ n4373) ) ;
 assign Ng26737 = ( (~ n3238) ) ;
 assign n3239 = ( Ng2165  &  (~ Ng2251) ) | ( (~ Ng2251)  &  n4375 ) | ( Ng2165  &  (~ n4375) ) ;
 assign Ng26736 = ( (~ n3239) ) ;
 assign n3240 = ( Ng2170  &  (~ Ng2247) ) | ( (~ Ng2247)  &  n4370 ) | ( Ng2170  &  (~ n4370) ) ;
 assign Ng26735 = ( (~ n3240) ) ;
 assign n3241 = ( (~ Ng2249)  &  Ng2170 ) | ( (~ Ng2249)  &  n4373 ) | ( Ng2170  &  (~ n4373) ) ;
 assign Ng26734 = ( (~ n3241) ) ;
 assign n3242 = ( Ng2170  &  (~ Ng2248) ) | ( (~ Ng2248)  &  n4375 ) | ( Ng2170  &  (~ n4375) ) ;
 assign Ng26733 = ( (~ n3242) ) ;
 assign n3243 = ( (~ Ng2244)  &  n4370 ) | ( (~ Ng2244)  &  n4385 ) | ( (~ n4370)  &  n4385 ) ;
 assign Ng26732 = ( (~ n3243) ) ;
 assign n3244 = ( (~ Ng2246)  &  n4373 ) | ( (~ Ng2246)  &  n4385 ) | ( (~ n4373)  &  n4385 ) ;
 assign Ng26731 = ( (~ n3244) ) ;
 assign n3245 = ( (~ Ng2245)  &  n4375 ) | ( (~ Ng2245)  &  n4385 ) | ( (~ n4375)  &  n4385 ) ;
 assign Ng26730 = ( (~ n3245) ) ;
 assign n3246 = ( (~ n763)  &  n765 ) | ( (~ n763)  &  (~ Ng2114) ) | ( (~ n765)  &  (~ Ng2114) ) ;
 assign Ng26728 = ( (~ n3246) ) ;
 assign n3247 = ( n760  &  (~ n763) ) | ( (~ n760)  &  (~ Ng2116) ) | ( (~ n763)  &  (~ Ng2116) ) ;
 assign Ng26727 = ( (~ n3247) ) ;
 assign n3248 = ( n754  &  (~ n763) ) | ( (~ n754)  &  (~ Ng2115) ) | ( (~ n763)  &  (~ Ng2115) ) ;
 assign Ng26726 = ( (~ n3248) ) ;
 assign n3249 = ( n1800  &  (~ Ng1559) ) | ( (~ Ng1559)  &  n4370 ) | ( n1800  &  (~ n4370) ) ;
 assign Ng26724 = ( (~ n3249) ) ;
 assign n3250 = ( n1800  &  (~ n4373) ) | ( n1800  &  (~ Ng1561) ) | ( n4373  &  (~ Ng1561) ) ;
 assign Ng26723 = ( (~ n3250) ) ;
 assign n3251 = ( n1800  &  (~ Ng1560) ) | ( (~ Ng1560)  &  n4375 ) | ( n1800  &  (~ n4375) ) ;
 assign Ng26722 = ( (~ n3251) ) ;
 assign n3252 = ( Ng1471  &  (~ Ng1556) ) | ( (~ Ng1556)  &  n4370 ) | ( Ng1471  &  (~ n4370) ) ;
 assign Ng26721 = ( (~ n3252) ) ;
 assign n3253 = ( (~ Ng1558)  &  Ng1471 ) | ( (~ Ng1558)  &  n4373 ) | ( Ng1471  &  (~ n4373) ) ;
 assign Ng26720 = ( (~ n3253) ) ;
 assign n3254 = ( Ng1471  &  (~ Ng1557) ) | ( (~ Ng1557)  &  n4375 ) | ( Ng1471  &  (~ n4375) ) ;
 assign Ng26719 = ( (~ n3254) ) ;
 assign n3255 = ( Ng1476  &  (~ Ng1553) ) | ( (~ Ng1553)  &  n4370 ) | ( Ng1476  &  (~ n4370) ) ;
 assign Ng26718 = ( (~ n3255) ) ;
 assign n3256 = ( (~ Ng1555)  &  Ng1476 ) | ( (~ Ng1555)  &  n4373 ) | ( Ng1476  &  (~ n4373) ) ;
 assign Ng26717 = ( (~ n3256) ) ;
 assign n3257 = ( Ng1476  &  (~ Ng1554) ) | ( (~ Ng1554)  &  n4375 ) | ( Ng1476  &  (~ n4375) ) ;
 assign Ng26716 = ( (~ n3257) ) ;
 assign n3258 = ( (~ Ng1550)  &  n4370 ) | ( (~ Ng1550)  &  n4404 ) | ( (~ n4370)  &  n4404 ) ;
 assign Ng26715 = ( (~ n3258) ) ;
 assign n3259 = ( (~ Ng1552)  &  n4373 ) | ( (~ Ng1552)  &  n4404 ) | ( (~ n4373)  &  n4404 ) ;
 assign Ng26714 = ( (~ n3259) ) ;
 assign n3260 = ( (~ Ng1551)  &  n4375 ) | ( (~ Ng1551)  &  n4404 ) | ( (~ n4375)  &  n4404 ) ;
 assign Ng26713 = ( (~ n3260) ) ;
 assign n3261 = ( (~ n756)  &  n758 ) | ( (~ n756)  &  (~ Ng1420) ) | ( (~ n758)  &  (~ Ng1420) ) ;
 assign Ng26711 = ( (~ n3261) ) ;
 assign n3262 = ( n753  &  (~ n756) ) | ( (~ n753)  &  (~ Ng1422) ) | ( (~ n756)  &  (~ Ng1422) ) ;
 assign Ng26710 = ( (~ n3262) ) ;
 assign n3263 = ( n747  &  (~ n756) ) | ( (~ n747)  &  (~ Ng1421) ) | ( (~ n756)  &  (~ Ng1421) ) ;
 assign Ng26709 = ( (~ n3263) ) ;
 assign n3264 = ( n1810  &  (~ Ng865) ) | ( (~ Ng865)  &  n4370 ) | ( n1810  &  (~ n4370) ) ;
 assign Ng26707 = ( (~ n3264) ) ;
 assign n3265 = ( n1810  &  (~ n4373) ) | ( n1810  &  (~ Ng867) ) | ( n4373  &  (~ Ng867) ) ;
 assign Ng26706 = ( (~ n3265) ) ;
 assign n3266 = ( n1810  &  (~ Ng866) ) | ( (~ Ng866)  &  n4375 ) | ( n1810  &  (~ n4375) ) ;
 assign Ng26705 = ( (~ n3266) ) ;
 assign n3267 = ( Ng785  &  (~ Ng862) ) | ( (~ Ng862)  &  n4370 ) | ( Ng785  &  (~ n4370) ) ;
 assign Ng26704 = ( (~ n3267) ) ;
 assign n3268 = ( (~ Ng864)  &  Ng785 ) | ( (~ Ng864)  &  n4373 ) | ( Ng785  &  (~ n4373) ) ;
 assign Ng26703 = ( (~ n3268) ) ;
 assign n3269 = ( Ng785  &  (~ Ng863) ) | ( (~ Ng863)  &  n4375 ) | ( Ng785  &  (~ n4375) ) ;
 assign Ng26702 = ( (~ n3269) ) ;
 assign n3270 = ( Ng789  &  (~ Ng859) ) | ( (~ Ng859)  &  n4370 ) | ( Ng789  &  (~ n4370) ) ;
 assign Ng26701 = ( (~ n3270) ) ;
 assign n3271 = ( (~ Ng861)  &  Ng789 ) | ( (~ Ng861)  &  n4373 ) | ( Ng789  &  (~ n4373) ) ;
 assign Ng26700 = ( (~ n3271) ) ;
 assign n3272 = ( Ng789  &  (~ Ng860) ) | ( (~ Ng860)  &  n4375 ) | ( Ng789  &  (~ n4375) ) ;
 assign Ng26699 = ( (~ n3272) ) ;
 assign n3273 = ( (~ Ng856)  &  n4370 ) | ( (~ Ng856)  &  n4423 ) | ( (~ n4370)  &  n4423 ) ;
 assign Ng26698 = ( (~ n3273) ) ;
 assign n3274 = ( (~ Ng858)  &  n4373 ) | ( (~ Ng858)  &  n4423 ) | ( (~ n4373)  &  n4423 ) ;
 assign Ng26697 = ( (~ n3274) ) ;
 assign n3275 = ( (~ Ng857)  &  n4375 ) | ( (~ Ng857)  &  n4423 ) | ( (~ n4375)  &  n4423 ) ;
 assign Ng26696 = ( (~ n3275) ) ;
 assign n3276 = ( (~ n749)  &  n751 ) | ( (~ n749)  &  (~ Ng734) ) | ( (~ n751)  &  (~ Ng734) ) ;
 assign Ng26694 = ( (~ n3276) ) ;
 assign n3277 = ( n746  &  (~ n749) ) | ( (~ n746)  &  (~ Ng736) ) | ( (~ n749)  &  (~ Ng736) ) ;
 assign Ng26693 = ( (~ n3277) ) ;
 assign n3278 = ( n743  &  (~ n749) ) | ( (~ n743)  &  (~ Ng735) ) | ( (~ n749)  &  (~ Ng735) ) ;
 assign Ng26692 = ( (~ n3278) ) ;
 assign n3279 = ( n1820  &  (~ Ng177) ) | ( (~ Ng177)  &  n4370 ) | ( n1820  &  (~ n4370) ) ;
 assign Ng26690 = ( (~ n3279) ) ;
 assign n3280 = ( n1820  &  (~ n4373) ) | ( n1820  &  (~ Ng179) ) | ( n4373  &  (~ Ng179) ) ;
 assign Ng26689 = ( (~ n3280) ) ;
 assign n3281 = ( n1820  &  (~ Ng178) ) | ( (~ Ng178)  &  n4375 ) | ( n1820  &  (~ n4375) ) ;
 assign Ng26688 = ( (~ n3281) ) ;
 assign n3282 = ( Ng97  &  (~ Ng174) ) | ( (~ Ng174)  &  n4370 ) | ( Ng97  &  (~ n4370) ) ;
 assign Ng26687 = ( (~ n3282) ) ;
 assign n3283 = ( (~ Ng176)  &  Ng97 ) | ( (~ Ng176)  &  n4373 ) | ( Ng97  &  (~ n4373) ) ;
 assign Ng26686 = ( (~ n3283) ) ;
 assign n3284 = ( Ng97  &  (~ Ng175) ) | ( (~ Ng175)  &  n4375 ) | ( Ng97  &  (~ n4375) ) ;
 assign Ng26685 = ( (~ n3284) ) ;
 assign n3285 = ( Ng101  &  (~ Ng171) ) | ( (~ Ng171)  &  n4370 ) | ( Ng101  &  (~ n4370) ) ;
 assign Ng26684 = ( (~ n3285) ) ;
 assign n3286 = ( Ng101  &  (~ Ng173) ) | ( (~ Ng173)  &  n4373 ) | ( Ng101  &  (~ n4373) ) ;
 assign Ng26683 = ( (~ n3286) ) ;
 assign n3287 = ( (~ Ng172)  &  Ng101 ) | ( (~ Ng172)  &  n4375 ) | ( Ng101  &  (~ n4375) ) ;
 assign Ng26682 = ( (~ n3287) ) ;
 assign n3288 = ( (~ Ng168)  &  n4370 ) | ( (~ Ng168)  &  n4442 ) | ( (~ n4370)  &  n4442 ) ;
 assign Ng26681 = ( (~ n3288) ) ;
 assign n3289 = ( (~ Ng170)  &  n4373 ) | ( (~ Ng170)  &  n4442 ) | ( (~ n4373)  &  n4442 ) ;
 assign Ng26680 = ( (~ n3289) ) ;
 assign n3290 = ( (~ Ng169)  &  n4375 ) | ( (~ Ng169)  &  n4442 ) | ( (~ n4375)  &  n4442 ) ;
 assign Ng26679 = ( (~ n3290) ) ;
 assign n3291 = ( (~ Ng1315)  &  (~ Ng2676) ) | ( Ng1315  &  n4445 ) | ( (~ Ng2676)  &  n4445 ) ;
 assign Ng26017 = ( (~ n3291) ) ;
 assign n3292 = ( (~ wire1603)  &  (~ Ng2673) ) | ( wire1603  &  n4445 ) | ( (~ Ng2673)  &  n4445 ) ;
 assign Ng26016 = ( (~ n3292) ) ;
 assign n3293 = ( (~ wire1605)  &  (~ Ng2670) ) | ( wire1605  &  n4445 ) | ( (~ Ng2670)  &  n4445 ) ;
 assign Ng26015 = ( (~ n3293) ) ;
 assign n3294 = ( (~ Ng1315)  &  (~ Ng2667) ) | ( Ng1315  &  n4446 ) | ( (~ Ng2667)  &  n4446 ) ;
 assign Ng26014 = ( (~ n3294) ) ;
 assign n3295 = ( (~ wire1603)  &  (~ Ng2664) ) | ( wire1603  &  n4446 ) | ( (~ Ng2664)  &  n4446 ) ;
 assign Ng26013 = ( (~ n3295) ) ;
 assign n3296 = ( (~ wire1605)  &  (~ Ng2661) ) | ( wire1605  &  n4446 ) | ( (~ Ng2661)  &  n4446 ) ;
 assign Ng26012 = ( (~ n3296) ) ;
 assign n3297 = ( Pg3229  &  Ng2366 ) | ( (~ Pg3229)  &  (~ Ng2380) ) | ( Ng2366  &  (~ Ng2380) ) ;
 assign Ng26011 = ( (~ n3297) ) ;
 assign n3298 = ( n1916  &  (~ Ng2160) ) | ( n1916  &  (~ n4447) ) | ( Ng2160  &  (~ n4447) ) ;
 assign Ng26010 = ( (~ n3298) ) ;
 assign n3299 = ( (~ Ng1315)  &  (~ Ng1982) ) | ( Ng1315  &  n4449 ) | ( (~ Ng1982)  &  n4449 ) ;
 assign Ng26008 = ( (~ n3299) ) ;
 assign n3300 = ( (~ wire1603)  &  (~ Ng1979) ) | ( wire1603  &  n4449 ) | ( (~ Ng1979)  &  n4449 ) ;
 assign Ng26007 = ( (~ n3300) ) ;
 assign n3301 = ( (~ wire1605)  &  (~ Ng1976) ) | ( wire1605  &  n4449 ) | ( (~ Ng1976)  &  n4449 ) ;
 assign Ng26006 = ( (~ n3301) ) ;
 assign n3302 = ( (~ Ng1315)  &  (~ Ng1973) ) | ( Ng1315  &  n4450 ) | ( (~ Ng1973)  &  n4450 ) ;
 assign Ng26005 = ( (~ n3302) ) ;
 assign n3303 = ( (~ wire1603)  &  (~ Ng1970) ) | ( wire1603  &  n4450 ) | ( (~ Ng1970)  &  n4450 ) ;
 assign Ng26004 = ( (~ n3303) ) ;
 assign n3304 = ( (~ wire1605)  &  (~ Ng1967) ) | ( wire1605  &  n4450 ) | ( (~ Ng1967)  &  n4450 ) ;
 assign Ng26003 = ( (~ n3304) ) ;
 assign n3305 = ( Pg3229  &  Ng1672 ) | ( (~ Pg3229)  &  (~ Ng1686) ) | ( Ng1672  &  (~ Ng1686) ) ;
 assign Ng26002 = ( (~ n3305) ) ;
 assign n3306 = ( n1916  &  (~ Ng1466) ) | ( n1916  &  (~ n4447) ) | ( Ng1466  &  (~ n4447) ) ;
 assign Ng26001 = ( (~ n3306) ) ;
 assign n3307 = ( (~ Ng1315)  &  (~ Ng1288) ) | ( Ng1315  &  n4451 ) | ( (~ Ng1288)  &  n4451 ) ;
 assign Ng25999 = ( (~ n3307) ) ;
 assign n3308 = ( (~ wire1603)  &  (~ Ng1285) ) | ( wire1603  &  n4451 ) | ( (~ Ng1285)  &  n4451 ) ;
 assign Ng25998 = ( (~ n3308) ) ;
 assign n3309 = ( (~ wire1605)  &  (~ Ng1282) ) | ( wire1605  &  n4451 ) | ( (~ Ng1282)  &  n4451 ) ;
 assign Ng25997 = ( (~ n3309) ) ;
 assign n3310 = ( (~ Ng1315)  &  (~ Ng1279) ) | ( Ng1315  &  n4452 ) | ( (~ Ng1279)  &  n4452 ) ;
 assign Ng25996 = ( (~ n3310) ) ;
 assign n3311 = ( (~ wire1603)  &  (~ Ng1276) ) | ( wire1603  &  n4452 ) | ( (~ Ng1276)  &  n4452 ) ;
 assign Ng25995 = ( (~ n3311) ) ;
 assign n3312 = ( (~ wire1605)  &  (~ Ng1273) ) | ( wire1605  &  n4452 ) | ( (~ Ng1273)  &  n4452 ) ;
 assign Ng25994 = ( (~ n3312) ) ;
 assign n3313 = ( Pg3229  &  Ng978 ) | ( (~ Pg3229)  &  (~ Ng992) ) | ( Ng978  &  (~ Ng992) ) ;
 assign Ng25993 = ( (~ n3313) ) ;
 assign n3314 = ( n1916  &  (~ Ng780) ) | ( n1916  &  (~ n4447) ) | ( Ng780  &  (~ n4447) ) ;
 assign Ng25992 = ( (~ n3314) ) ;
 assign n3315 = ( (~ Ng1315)  &  (~ Ng602) ) | ( Ng1315  &  n4453 ) | ( (~ Ng602)  &  n4453 ) ;
 assign Ng25990 = ( (~ n3315) ) ;
 assign n3316 = ( (~ wire1603)  &  (~ Ng599) ) | ( wire1603  &  n4453 ) | ( (~ Ng599)  &  n4453 ) ;
 assign Ng25989 = ( (~ n3316) ) ;
 assign n3317 = ( (~ wire1605)  &  (~ Ng596) ) | ( wire1605  &  n4453 ) | ( (~ Ng596)  &  n4453 ) ;
 assign Ng25988 = ( (~ n3317) ) ;
 assign n3318 = ( (~ Ng1315)  &  (~ Ng593) ) | ( Ng1315  &  n4454 ) | ( (~ Ng593)  &  n4454 ) ;
 assign Ng25987 = ( (~ n3318) ) ;
 assign n3319 = ( (~ wire1603)  &  (~ Ng590) ) | ( wire1603  &  n4454 ) | ( (~ Ng590)  &  n4454 ) ;
 assign Ng25986 = ( (~ n3319) ) ;
 assign n3320 = ( (~ wire1605)  &  (~ Ng587) ) | ( wire1605  &  n4454 ) | ( (~ Ng587)  &  n4454 ) ;
 assign Ng25985 = ( (~ n3320) ) ;
 assign n3321 = ( Pg3229  &  Ng291 ) | ( (~ Pg3229)  &  (~ Ng305) ) | ( Ng291  &  (~ Ng305) ) ;
 assign Ng25984 = ( (~ n3321) ) ;
 assign n3322 = ( n1916  &  (~ Ng92) ) | ( n1916  &  (~ n4447) ) | ( Ng92  &  (~ n4447) ) ;
 assign Ng25983 = ( (~ n3322) ) ;
 assign n3323 = ( (~ Ng3147)  &  (~ n4455) ) | ( n2503  &  (~ n4455) ) | ( (~ Ng3097)  &  (~ n4455) ) ;
 assign n3324 = ( wire1612  &  n733 ) | ( (~ wire1612)  &  (~ Ng11593) ) | ( n733  &  (~ Ng11593) ) ;
 assign Ng25172 = ( (~ n3324) ) ;
 assign n3325 = ( Ng853  &  n1546 ) | ( (~ Ng853)  &  (~ Ng2554) ) | ( n1546  &  (~ Ng2554) ) ;
 assign Ng25171 = ( (~ n3325) ) ;
 assign n3326 = ( (~ wire1594)  &  (~ Ng2553) ) | ( wire1594  &  n1546 ) | ( (~ Ng2553)  &  n1546 ) ;
 assign Ng25170 = ( (~ n3326) ) ;
 assign n3327 = ( wire1612  &  n1546 ) | ( (~ wire1612)  &  (~ Ng2552) ) | ( n1546  &  (~ Ng2552) ) ;
 assign Ng25169 = ( (~ n3327) ) ;
 assign n3328 = ( Ng853  &  n1889 ) | ( (~ Ng853)  &  (~ Ng11595) ) | ( n1889  &  (~ Ng11595) ) ;
 assign Ng25168 = ( (~ n3328) ) ;
 assign n3329 = ( wire1594  &  n1889 ) | ( (~ wire1594)  &  (~ Ng11594) ) | ( n1889  &  (~ Ng11594) ) ;
 assign Ng25167 = ( (~ n3329) ) ;
 assign n3330 = ( wire1612  &  n1889 ) | ( (~ wire1612)  &  (~ Ng11598) ) | ( n1889  &  (~ Ng11598) ) ;
 assign Ng25166 = ( (~ n3330) ) ;
 assign n3331 = ( Ng853  &  n733 ) | ( (~ Ng853)  &  (~ Ng11597) ) | ( n733  &  (~ Ng11597) ) ;
 assign Ng25165 = ( (~ n3331) ) ;
 assign n3332 = ( wire1594  &  n733 ) | ( (~ wire1594)  &  (~ Ng11596) ) | ( n733  &  (~ Ng11596) ) ;
 assign Ng25164 = ( (~ n3332) ) ;
 assign n3333 = ( wire1612  &  n730 ) | ( (~ wire1612)  &  (~ Ng11566) ) | ( n730  &  (~ Ng11566) ) ;
 assign Ng25161 = ( (~ n3333) ) ;
 assign n3334 = ( Ng853  &  n1556 ) | ( (~ Ng853)  &  (~ Ng1860) ) | ( n1556  &  (~ Ng1860) ) ;
 assign Ng25160 = ( (~ n3334) ) ;
 assign n3335 = ( (~ wire1594)  &  (~ Ng1859) ) | ( wire1594  &  n1556 ) | ( (~ Ng1859)  &  n1556 ) ;
 assign Ng25159 = ( (~ n3335) ) ;
 assign n3336 = ( wire1612  &  n1556 ) | ( (~ wire1612)  &  (~ Ng1858) ) | ( n1556  &  (~ Ng1858) ) ;
 assign Ng25158 = ( (~ n3336) ) ;
 assign n3337 = ( Ng853  &  n1893 ) | ( (~ Ng853)  &  (~ Ng11568) ) | ( n1893  &  (~ Ng11568) ) ;
 assign Ng25157 = ( (~ n3337) ) ;
 assign n3338 = ( wire1594  &  n1893 ) | ( (~ wire1594)  &  (~ Ng11567) ) | ( n1893  &  (~ Ng11567) ) ;
 assign Ng25156 = ( (~ n3338) ) ;
 assign n3339 = ( wire1612  &  n1893 ) | ( (~ wire1612)  &  (~ Ng11571) ) | ( n1893  &  (~ Ng11571) ) ;
 assign Ng25155 = ( (~ n3339) ) ;
 assign n3340 = ( Ng853  &  n730 ) | ( (~ Ng853)  &  (~ Ng11570) ) | ( n730  &  (~ Ng11570) ) ;
 assign Ng25154 = ( (~ n3340) ) ;
 assign n3341 = ( wire1594  &  n730 ) | ( (~ wire1594)  &  (~ Ng11569) ) | ( n730  &  (~ Ng11569) ) ;
 assign Ng25153 = ( (~ n3341) ) ;
 assign n3342 = ( wire1612  &  n726 ) | ( (~ wire1612)  &  (~ Ng11539) ) | ( n726  &  (~ Ng11539) ) ;
 assign Ng25150 = ( (~ n3342) ) ;
 assign n3343 = ( Ng853  &  n1566 ) | ( (~ Ng853)  &  (~ Ng1166) ) | ( n1566  &  (~ Ng1166) ) ;
 assign Ng25149 = ( (~ n3343) ) ;
 assign n3344 = ( (~ wire1594)  &  (~ Ng1165) ) | ( wire1594  &  n1566 ) | ( (~ Ng1165)  &  n1566 ) ;
 assign Ng25148 = ( (~ n3344) ) ;
 assign n3345 = ( wire1612  &  n1566 ) | ( (~ wire1612)  &  (~ Ng1164) ) | ( n1566  &  (~ Ng1164) ) ;
 assign Ng25147 = ( (~ n3345) ) ;
 assign n3346 = ( Ng853  &  n1897 ) | ( (~ Ng853)  &  (~ Ng11541) ) | ( n1897  &  (~ Ng11541) ) ;
 assign Ng25146 = ( (~ n3346) ) ;
 assign n3347 = ( wire1594  &  n1897 ) | ( (~ wire1594)  &  (~ Ng11540) ) | ( n1897  &  (~ Ng11540) ) ;
 assign Ng25145 = ( (~ n3347) ) ;
 assign n3348 = ( wire1612  &  n1897 ) | ( (~ wire1612)  &  (~ Ng11544) ) | ( n1897  &  (~ Ng11544) ) ;
 assign Ng25144 = ( (~ n3348) ) ;
 assign n3349 = ( Ng853  &  n726 ) | ( (~ Ng853)  &  (~ Ng11543) ) | ( n726  &  (~ Ng11543) ) ;
 assign Ng25143 = ( (~ n3349) ) ;
 assign n3350 = ( wire1594  &  n726 ) | ( (~ wire1594)  &  (~ Ng11542) ) | ( n726  &  (~ Ng11542) ) ;
 assign Ng25142 = ( (~ n3350) ) ;
 assign n3351 = ( wire1612  &  n722 ) | ( (~ wire1612)  &  (~ Ng11512) ) | ( n722  &  (~ Ng11512) ) ;
 assign Ng25139 = ( (~ n3351) ) ;
 assign n3352 = ( Ng853  &  n1576 ) | ( (~ Ng853)  &  (~ Ng479) ) | ( n1576  &  (~ Ng479) ) ;
 assign Ng25138 = ( (~ n3352) ) ;
 assign n3353 = ( (~ wire1594)  &  (~ Ng478) ) | ( wire1594  &  n1576 ) | ( (~ Ng478)  &  n1576 ) ;
 assign Ng25137 = ( (~ n3353) ) ;
 assign n3354 = ( wire1612  &  n1576 ) | ( (~ wire1612)  &  (~ Ng477) ) | ( n1576  &  (~ Ng477) ) ;
 assign Ng25136 = ( (~ n3354) ) ;
 assign n3355 = ( Ng853  &  n1901 ) | ( (~ Ng853)  &  (~ Ng11514) ) | ( n1901  &  (~ Ng11514) ) ;
 assign Ng25135 = ( (~ n3355) ) ;
 assign n3356 = ( wire1594  &  n1901 ) | ( (~ wire1594)  &  (~ Ng11513) ) | ( n1901  &  (~ Ng11513) ) ;
 assign Ng25134 = ( (~ n3356) ) ;
 assign n3357 = ( wire1612  &  n1901 ) | ( (~ wire1612)  &  (~ Ng11517) ) | ( n1901  &  (~ Ng11517) ) ;
 assign Ng25133 = ( (~ n3357) ) ;
 assign n3358 = ( Ng853  &  n722 ) | ( (~ Ng853)  &  (~ Ng11516) ) | ( n722  &  (~ Ng11516) ) ;
 assign Ng25132 = ( (~ n3358) ) ;
 assign n3359 = ( wire1594  &  n722 ) | ( (~ wire1594)  &  (~ Ng11515) ) | ( n722  &  (~ Ng11515) ) ;
 assign Ng25131 = ( (~ n3359) ) ;
 assign n3360 = ( Ng853  &  n488 ) | ( (~ Ng853)  &  (~ Ng2563) ) | ( n488  &  (~ Ng2563) ) ;
 assign Ng24417 = ( (~ n3360) ) ;
 assign n3361 = ( (~ wire1594)  &  (~ Ng2562) ) | ( wire1594  &  n488 ) | ( (~ Ng2562)  &  n488 ) ;
 assign Ng24416 = ( (~ n3361) ) ;
 assign n3362 = ( wire1612  &  n488 ) | ( (~ wire1612)  &  (~ Ng2561) ) | ( n488  &  (~ Ng2561) ) ;
 assign Ng24415 = ( (~ n3362) ) ;
 assign n3363 = ( Ng853  &  (~ n629) ) | ( (~ Ng853)  &  (~ Ng2539) ) | ( (~ n629)  &  (~ Ng2539) ) ;
 assign Ng24414 = ( (~ n3363) ) ;
 assign n3364 = ( (~ wire1594)  &  (~ Ng2559) ) | ( wire1594  &  (~ n629) ) | ( (~ Ng2559)  &  (~ n629) ) ;
 assign Ng24413 = ( (~ n3364) ) ;
 assign n3365 = ( wire1612  &  (~ n629) ) | ( (~ wire1612)  &  (~ Ng2555) ) | ( (~ n629)  &  (~ Ng2555) ) ;
 assign Ng24412 = ( (~ n3365) ) ;
 assign n3366 = ( (~ n640)  &  (~ n2450) ) | ( (~ n640)  &  (~ Ng2238) ) | ( n2450  &  (~ Ng2238) ) ;
 assign Ng24411 = ( (~ n3366) ) ;
 assign n3367 = ( (~ Ng2240)  &  (~ n640) ) | ( (~ Ng2240)  &  n4503 ) | ( (~ n640)  &  (~ n4503) ) ;
 assign Ng24410 = ( (~ n3367) ) ;
 assign n3368 = ( (~ n640)  &  (~ Ng2239) ) | ( (~ Ng2239)  &  n4506 ) | ( (~ n640)  &  (~ n4506) ) ;
 assign Ng24409 = ( (~ n3368) ) ;
 assign n3369 = ( (~ n642)  &  (~ n2450) ) | ( (~ n642)  &  (~ Ng2235) ) | ( n2450  &  (~ Ng2235) ) ;
 assign Ng24408 = ( (~ n3369) ) ;
 assign n3370 = ( (~ Ng2237)  &  (~ n642) ) | ( (~ Ng2237)  &  n4503 ) | ( (~ n642)  &  (~ n4503) ) ;
 assign Ng24407 = ( (~ n3370) ) ;
 assign n3371 = ( (~ n642)  &  (~ Ng2236) ) | ( (~ Ng2236)  &  n4506 ) | ( (~ n642)  &  (~ n4506) ) ;
 assign Ng24406 = ( (~ n3371) ) ;
 assign n3372 = ( Ng2200  &  (~ n2450) ) | ( Ng2200  &  (~ Ng2232) ) | ( n2450  &  (~ Ng2232) ) ;
 assign Ng24405 = ( (~ n3372) ) ;
 assign n3373 = ( (~ Ng2234)  &  Ng2200 ) | ( (~ Ng2234)  &  n4503 ) | ( Ng2200  &  (~ n4503) ) ;
 assign Ng24404 = ( (~ n3373) ) ;
 assign n3374 = ( Ng2200  &  (~ Ng2233) ) | ( (~ Ng2233)  &  n4506 ) | ( Ng2200  &  (~ n4506) ) ;
 assign Ng24403 = ( (~ n3374) ) ;
 assign n3375 = ( Ng2195  &  (~ n2450) ) | ( Ng2195  &  (~ Ng2229) ) | ( n2450  &  (~ Ng2229) ) ;
 assign Ng24402 = ( (~ n3375) ) ;
 assign n3376 = ( (~ Ng2231)  &  Ng2195 ) | ( (~ Ng2231)  &  n4503 ) | ( Ng2195  &  (~ n4503) ) ;
 assign Ng24401 = ( (~ n3376) ) ;
 assign n3377 = ( Ng2195  &  (~ Ng2230) ) | ( (~ Ng2230)  &  n4506 ) | ( Ng2195  &  (~ n4506) ) ;
 assign Ng24400 = ( (~ n3377) ) ;
 assign n3378 = ( Ng2190  &  (~ n2450) ) | ( Ng2190  &  (~ Ng2226) ) | ( n2450  &  (~ Ng2226) ) ;
 assign Ng24399 = ( (~ n3378) ) ;
 assign n3379 = ( (~ Ng2228)  &  Ng2190 ) | ( (~ Ng2228)  &  n4503 ) | ( Ng2190  &  (~ n4503) ) ;
 assign Ng24398 = ( (~ n3379) ) ;
 assign n3380 = ( Ng2190  &  (~ Ng2227) ) | ( (~ Ng2227)  &  n4506 ) | ( Ng2190  &  (~ n4506) ) ;
 assign Ng24397 = ( (~ n3380) ) ;
 assign n3381 = ( Ng2185  &  (~ n2450) ) | ( Ng2185  &  (~ Ng2223) ) | ( n2450  &  (~ Ng2223) ) ;
 assign Ng24396 = ( (~ n3381) ) ;
 assign n3382 = ( (~ Ng2225)  &  Ng2185 ) | ( (~ Ng2225)  &  n4503 ) | ( Ng2185  &  (~ n4503) ) ;
 assign Ng24395 = ( (~ n3382) ) ;
 assign n3383 = ( Ng2185  &  (~ Ng2224) ) | ( (~ Ng2224)  &  n4506 ) | ( Ng2185  &  (~ n4506) ) ;
 assign Ng24394 = ( (~ n3383) ) ;
 assign n3384 = ( Ng2180  &  (~ n2450) ) | ( Ng2180  &  (~ Ng2220) ) | ( n2450  &  (~ Ng2220) ) ;
 assign Ng24393 = ( (~ n3384) ) ;
 assign n3385 = ( (~ Ng2222)  &  Ng2180 ) | ( (~ Ng2222)  &  n4503 ) | ( Ng2180  &  (~ n4503) ) ;
 assign Ng24392 = ( (~ n3385) ) ;
 assign n3386 = ( Ng2180  &  (~ Ng2221) ) | ( (~ Ng2221)  &  n4506 ) | ( Ng2180  &  (~ n4506) ) ;
 assign Ng24391 = ( (~ n3386) ) ;
 assign n3387 = ( Ng2175  &  (~ n2450) ) | ( Ng2175  &  (~ Ng2217) ) | ( n2450  &  (~ Ng2217) ) ;
 assign Ng24390 = ( (~ n3387) ) ;
 assign n3388 = ( Ng2175  &  (~ Ng2219) ) | ( (~ Ng2219)  &  n4503 ) | ( Ng2175  &  (~ n4503) ) ;
 assign Ng24389 = ( (~ n3388) ) ;
 assign n3389 = ( (~ Ng2218)  &  Ng2175 ) | ( (~ Ng2218)  &  n4506 ) | ( Ng2175  &  (~ n4506) ) ;
 assign Ng24388 = ( (~ n3389) ) ;
 assign n3390 = ( Ng2170  &  (~ n2450) ) | ( Ng2170  &  (~ Ng2208) ) | ( n2450  &  (~ Ng2208) ) ;
 assign Ng24387 = ( (~ n3390) ) ;
 assign n3391 = ( (~ Ng2210)  &  Ng2170 ) | ( (~ Ng2210)  &  n4503 ) | ( Ng2170  &  (~ n4503) ) ;
 assign Ng24386 = ( (~ n3391) ) ;
 assign n3392 = ( Ng2170  &  (~ Ng2209) ) | ( (~ Ng2209)  &  n4506 ) | ( Ng2170  &  (~ n4506) ) ;
 assign Ng24385 = ( (~ n3392) ) ;
 assign n3393 = ( Ng2165  &  (~ n2450) ) | ( Ng2165  &  (~ Ng2205) ) | ( n2450  &  (~ Ng2205) ) ;
 assign Ng24384 = ( (~ n3393) ) ;
 assign n3394 = ( (~ Ng2207)  &  Ng2165 ) | ( (~ Ng2207)  &  n4503 ) | ( Ng2165  &  (~ n4503) ) ;
 assign Ng24383 = ( (~ n3394) ) ;
 assign n3395 = ( Ng2165  &  (~ Ng2206) ) | ( (~ Ng2206)  &  n4506 ) | ( Ng2165  &  (~ n4506) ) ;
 assign Ng24382 = ( (~ n3395) ) ;
 assign n3396 = ( Ng853  &  n443 ) | ( (~ Ng853)  &  (~ Ng1869) ) | ( n443  &  (~ Ng1869) ) ;
 assign Ng24376 = ( (~ n3396) ) ;
 assign n3397 = ( (~ wire1594)  &  (~ Ng1868) ) | ( wire1594  &  n443 ) | ( (~ Ng1868)  &  n443 ) ;
 assign Ng24375 = ( (~ n3397) ) ;
 assign n3398 = ( wire1612  &  n443 ) | ( (~ wire1612)  &  (~ Ng1867) ) | ( n443  &  (~ Ng1867) ) ;
 assign Ng24374 = ( (~ n3398) ) ;
 assign n3399 = ( Ng853  &  (~ n615) ) | ( (~ Ng853)  &  (~ Ng1845) ) | ( (~ n615)  &  (~ Ng1845) ) ;
 assign Ng24373 = ( (~ n3399) ) ;
 assign n3400 = ( (~ wire1594)  &  (~ Ng1865) ) | ( wire1594  &  (~ n615) ) | ( (~ Ng1865)  &  (~ n615) ) ;
 assign Ng24372 = ( (~ n3400) ) ;
 assign n3401 = ( wire1612  &  (~ n615) ) | ( (~ wire1612)  &  (~ Ng1861) ) | ( (~ n615)  &  (~ Ng1861) ) ;
 assign Ng24371 = ( (~ n3401) ) ;
 assign n3402 = ( (~ n636)  &  (~ n2450) ) | ( (~ n636)  &  (~ Ng1544) ) | ( n2450  &  (~ Ng1544) ) ;
 assign Ng24370 = ( (~ n3402) ) ;
 assign n3403 = ( (~ Ng1546)  &  (~ n636) ) | ( (~ Ng1546)  &  n4503 ) | ( (~ n636)  &  (~ n4503) ) ;
 assign Ng24369 = ( (~ n3403) ) ;
 assign n3404 = ( (~ n636)  &  (~ Ng1545) ) | ( (~ Ng1545)  &  n4506 ) | ( (~ n636)  &  (~ n4506) ) ;
 assign Ng24368 = ( (~ n3404) ) ;
 assign n3405 = ( (~ n638)  &  (~ n2450) ) | ( (~ n638)  &  (~ Ng1541) ) | ( n2450  &  (~ Ng1541) ) ;
 assign Ng24367 = ( (~ n3405) ) ;
 assign n3406 = ( (~ Ng1543)  &  (~ n638) ) | ( (~ Ng1543)  &  n4503 ) | ( (~ n638)  &  (~ n4503) ) ;
 assign Ng24366 = ( (~ n3406) ) ;
 assign n3407 = ( (~ n638)  &  (~ Ng1542) ) | ( (~ Ng1542)  &  n4506 ) | ( (~ n638)  &  (~ n4506) ) ;
 assign Ng24365 = ( (~ n3407) ) ;
 assign n3408 = ( Ng1506  &  (~ n2450) ) | ( Ng1506  &  (~ Ng1538) ) | ( n2450  &  (~ Ng1538) ) ;
 assign Ng24364 = ( (~ n3408) ) ;
 assign n3409 = ( (~ Ng1540)  &  Ng1506 ) | ( (~ Ng1540)  &  n4503 ) | ( Ng1506  &  (~ n4503) ) ;
 assign Ng24363 = ( (~ n3409) ) ;
 assign n3410 = ( Ng1506  &  (~ Ng1539) ) | ( (~ Ng1539)  &  n4506 ) | ( Ng1506  &  (~ n4506) ) ;
 assign Ng24362 = ( (~ n3410) ) ;
 assign n3411 = ( Ng1501  &  (~ n2450) ) | ( Ng1501  &  (~ Ng1535) ) | ( n2450  &  (~ Ng1535) ) ;
 assign Ng24361 = ( (~ n3411) ) ;
 assign n3412 = ( (~ Ng1537)  &  Ng1501 ) | ( (~ Ng1537)  &  n4503 ) | ( Ng1501  &  (~ n4503) ) ;
 assign Ng24360 = ( (~ n3412) ) ;
 assign n3413 = ( Ng1501  &  (~ Ng1536) ) | ( (~ Ng1536)  &  n4506 ) | ( Ng1501  &  (~ n4506) ) ;
 assign Ng24359 = ( (~ n3413) ) ;
 assign n3414 = ( Ng1496  &  (~ n2450) ) | ( Ng1496  &  (~ Ng1532) ) | ( n2450  &  (~ Ng1532) ) ;
 assign Ng24358 = ( (~ n3414) ) ;
 assign n3415 = ( (~ Ng1534)  &  Ng1496 ) | ( (~ Ng1534)  &  n4503 ) | ( Ng1496  &  (~ n4503) ) ;
 assign Ng24357 = ( (~ n3415) ) ;
 assign n3416 = ( Ng1496  &  (~ Ng1533) ) | ( (~ Ng1533)  &  n4506 ) | ( Ng1496  &  (~ n4506) ) ;
 assign Ng24356 = ( (~ n3416) ) ;
 assign n3417 = ( Ng1491  &  (~ n2450) ) | ( Ng1491  &  (~ Ng1529) ) | ( n2450  &  (~ Ng1529) ) ;
 assign Ng24355 = ( (~ n3417) ) ;
 assign n3418 = ( (~ Ng1531)  &  Ng1491 ) | ( (~ Ng1531)  &  n4503 ) | ( Ng1491  &  (~ n4503) ) ;
 assign Ng24354 = ( (~ n3418) ) ;
 assign n3419 = ( Ng1491  &  (~ Ng1530) ) | ( (~ Ng1530)  &  n4506 ) | ( Ng1491  &  (~ n4506) ) ;
 assign Ng24353 = ( (~ n3419) ) ;
 assign n3420 = ( Ng1486  &  (~ n2450) ) | ( Ng1486  &  (~ Ng1526) ) | ( n2450  &  (~ Ng1526) ) ;
 assign Ng24352 = ( (~ n3420) ) ;
 assign n3421 = ( Ng1486  &  (~ Ng1528) ) | ( (~ Ng1528)  &  n4503 ) | ( Ng1486  &  (~ n4503) ) ;
 assign Ng24351 = ( (~ n3421) ) ;
 assign n3422 = ( (~ Ng1527)  &  Ng1486 ) | ( (~ Ng1527)  &  n4506 ) | ( Ng1486  &  (~ n4506) ) ;
 assign Ng24350 = ( (~ n3422) ) ;
 assign n3423 = ( Ng1481  &  (~ n2450) ) | ( Ng1481  &  (~ Ng1523) ) | ( n2450  &  (~ Ng1523) ) ;
 assign Ng24349 = ( (~ n3423) ) ;
 assign n3424 = ( Ng1481  &  (~ Ng1525) ) | ( (~ Ng1525)  &  n4503 ) | ( Ng1481  &  (~ n4503) ) ;
 assign Ng24348 = ( (~ n3424) ) ;
 assign n3425 = ( (~ Ng1524)  &  Ng1481 ) | ( (~ Ng1524)  &  n4506 ) | ( Ng1481  &  (~ n4506) ) ;
 assign Ng24347 = ( (~ n3425) ) ;
 assign n3426 = ( Ng1476  &  (~ n2450) ) | ( Ng1476  &  (~ Ng1514) ) | ( n2450  &  (~ Ng1514) ) ;
 assign Ng24346 = ( (~ n3426) ) ;
 assign n3427 = ( (~ Ng1516)  &  Ng1476 ) | ( (~ Ng1516)  &  n4503 ) | ( Ng1476  &  (~ n4503) ) ;
 assign Ng24345 = ( (~ n3427) ) ;
 assign n3428 = ( Ng1476  &  (~ Ng1515) ) | ( (~ Ng1515)  &  n4506 ) | ( Ng1476  &  (~ n4506) ) ;
 assign Ng24344 = ( (~ n3428) ) ;
 assign n3429 = ( Ng1471  &  (~ n2450) ) | ( Ng1471  &  (~ Ng1511) ) | ( n2450  &  (~ Ng1511) ) ;
 assign Ng24343 = ( (~ n3429) ) ;
 assign n3430 = ( (~ Ng1513)  &  Ng1471 ) | ( (~ Ng1513)  &  n4503 ) | ( Ng1471  &  (~ n4503) ) ;
 assign Ng24342 = ( (~ n3430) ) ;
 assign n3431 = ( Ng1471  &  (~ Ng1512) ) | ( (~ Ng1512)  &  n4506 ) | ( Ng1471  &  (~ n4506) ) ;
 assign Ng24341 = ( (~ n3431) ) ;
 assign n3432 = ( Ng853  &  n393 ) | ( (~ Ng853)  &  (~ Ng1175) ) | ( n393  &  (~ Ng1175) ) ;
 assign Ng24335 = ( (~ n3432) ) ;
 assign n3433 = ( (~ wire1594)  &  (~ Ng1174) ) | ( wire1594  &  n393 ) | ( (~ Ng1174)  &  n393 ) ;
 assign Ng24334 = ( (~ n3433) ) ;
 assign n3434 = ( wire1612  &  n393 ) | ( (~ wire1612)  &  (~ Ng1173) ) | ( n393  &  (~ Ng1173) ) ;
 assign Ng24333 = ( (~ n3434) ) ;
 assign n3435 = ( Ng853  &  (~ n601) ) | ( (~ Ng853)  &  (~ Ng1151) ) | ( (~ n601)  &  (~ Ng1151) ) ;
 assign Ng24332 = ( (~ n3435) ) ;
 assign n3436 = ( (~ wire1594)  &  (~ Ng1171) ) | ( wire1594  &  (~ n601) ) | ( (~ Ng1171)  &  (~ n601) ) ;
 assign Ng24331 = ( (~ n3436) ) ;
 assign n3437 = ( wire1612  &  (~ n601) ) | ( (~ wire1612)  &  (~ Ng1167) ) | ( (~ n601)  &  (~ Ng1167) ) ;
 assign Ng24330 = ( (~ n3437) ) ;
 assign n3438 = ( (~ n627)  &  (~ n2450) ) | ( (~ n627)  &  (~ Ng850) ) | ( n2450  &  (~ Ng850) ) ;
 assign Ng24329 = ( (~ n3438) ) ;
 assign n3439 = ( (~ Ng852)  &  (~ n627) ) | ( (~ Ng852)  &  n4503 ) | ( (~ n627)  &  (~ n4503) ) ;
 assign Ng24328 = ( (~ n3439) ) ;
 assign n3440 = ( (~ n627)  &  (~ Ng851) ) | ( (~ Ng851)  &  n4506 ) | ( (~ n627)  &  (~ n4506) ) ;
 assign Ng24327 = ( (~ n3440) ) ;
 assign n3441 = ( (~ n634)  &  (~ n2450) ) | ( (~ n634)  &  (~ Ng847) ) | ( n2450  &  (~ Ng847) ) ;
 assign Ng24326 = ( (~ n3441) ) ;
 assign n3442 = ( (~ Ng849)  &  (~ n634) ) | ( (~ Ng849)  &  n4503 ) | ( (~ n634)  &  (~ n4503) ) ;
 assign Ng24325 = ( (~ n3442) ) ;
 assign n3443 = ( (~ n634)  &  (~ Ng848) ) | ( (~ Ng848)  &  n4506 ) | ( (~ n634)  &  (~ n4506) ) ;
 assign Ng24324 = ( (~ n3443) ) ;
 assign n3444 = ( Ng813  &  (~ n2450) ) | ( Ng813  &  (~ Ng844) ) | ( n2450  &  (~ Ng844) ) ;
 assign Ng24323 = ( (~ n3444) ) ;
 assign n3445 = ( (~ Ng846)  &  Ng813 ) | ( (~ Ng846)  &  n4503 ) | ( Ng813  &  (~ n4503) ) ;
 assign Ng24322 = ( (~ n3445) ) ;
 assign n3446 = ( Ng813  &  (~ Ng845) ) | ( (~ Ng845)  &  n4506 ) | ( Ng813  &  (~ n4506) ) ;
 assign Ng24321 = ( (~ n3446) ) ;
 assign n3447 = ( Ng809  &  (~ n2450) ) | ( Ng809  &  (~ Ng841) ) | ( n2450  &  (~ Ng841) ) ;
 assign Ng24320 = ( (~ n3447) ) ;
 assign n3448 = ( (~ Ng843)  &  Ng809 ) | ( (~ Ng843)  &  n4503 ) | ( Ng809  &  (~ n4503) ) ;
 assign Ng24319 = ( (~ n3448) ) ;
 assign n3449 = ( Ng809  &  (~ Ng842) ) | ( (~ Ng842)  &  n4506 ) | ( Ng809  &  (~ n4506) ) ;
 assign Ng24318 = ( (~ n3449) ) ;
 assign n3450 = ( Ng805  &  (~ n2450) ) | ( Ng805  &  (~ Ng838) ) | ( n2450  &  (~ Ng838) ) ;
 assign Ng24317 = ( (~ n3450) ) ;
 assign n3451 = ( (~ Ng840)  &  Ng805 ) | ( (~ Ng840)  &  n4503 ) | ( Ng805  &  (~ n4503) ) ;
 assign Ng24316 = ( (~ n3451) ) ;
 assign n3452 = ( Ng805  &  (~ Ng839) ) | ( (~ Ng839)  &  n4506 ) | ( Ng805  &  (~ n4506) ) ;
 assign Ng24315 = ( (~ n3452) ) ;
 assign n3453 = ( Ng801  &  (~ n2450) ) | ( Ng801  &  (~ Ng835) ) | ( n2450  &  (~ Ng835) ) ;
 assign Ng24314 = ( (~ n3453) ) ;
 assign n3454 = ( Ng801  &  (~ Ng837) ) | ( (~ Ng837)  &  n4503 ) | ( Ng801  &  (~ n4503) ) ;
 assign Ng24313 = ( (~ n3454) ) ;
 assign n3455 = ( (~ Ng836)  &  Ng801 ) | ( (~ Ng836)  &  n4506 ) | ( Ng801  &  (~ n4506) ) ;
 assign Ng24312 = ( (~ n3455) ) ;
 assign n3456 = ( Ng797  &  (~ n2450) ) | ( Ng797  &  (~ Ng832) ) | ( n2450  &  (~ Ng832) ) ;
 assign Ng24311 = ( (~ n3456) ) ;
 assign n3457 = ( Ng797  &  (~ Ng834) ) | ( (~ Ng834)  &  n4503 ) | ( Ng797  &  (~ n4503) ) ;
 assign Ng24310 = ( (~ n3457) ) ;
 assign n3458 = ( (~ Ng833)  &  Ng797 ) | ( (~ Ng833)  &  n4506 ) | ( Ng797  &  (~ n4506) ) ;
 assign Ng24309 = ( (~ n3458) ) ;
 assign n3459 = ( Ng793  &  (~ n2450) ) | ( Ng793  &  (~ Ng829) ) | ( n2450  &  (~ Ng829) ) ;
 assign Ng24308 = ( (~ n3459) ) ;
 assign n3460 = ( Ng793  &  (~ Ng831) ) | ( (~ Ng831)  &  n4503 ) | ( Ng793  &  (~ n4503) ) ;
 assign Ng24307 = ( (~ n3460) ) ;
 assign n3461 = ( (~ Ng830)  &  Ng793 ) | ( (~ Ng830)  &  n4506 ) | ( Ng793  &  (~ n4506) ) ;
 assign Ng24306 = ( (~ n3461) ) ;
 assign n3462 = ( Ng789  &  (~ n2450) ) | ( Ng789  &  (~ Ng820) ) | ( n2450  &  (~ Ng820) ) ;
 assign Ng24305 = ( (~ n3462) ) ;
 assign n3463 = ( (~ Ng822)  &  Ng789 ) | ( (~ Ng822)  &  n4503 ) | ( Ng789  &  (~ n4503) ) ;
 assign Ng24304 = ( (~ n3463) ) ;
 assign n3464 = ( Ng789  &  (~ Ng821) ) | ( (~ Ng821)  &  n4506 ) | ( Ng789  &  (~ n4506) ) ;
 assign Ng24303 = ( (~ n3464) ) ;
 assign n3465 = ( Ng785  &  (~ n2450) ) | ( Ng785  &  (~ Ng817) ) | ( n2450  &  (~ Ng817) ) ;
 assign Ng24302 = ( (~ n3465) ) ;
 assign n3466 = ( (~ Ng819)  &  Ng785 ) | ( (~ Ng819)  &  n4503 ) | ( Ng785  &  (~ n4503) ) ;
 assign Ng24301 = ( (~ n3466) ) ;
 assign n3467 = ( Ng785  &  (~ Ng818) ) | ( (~ Ng818)  &  n4506 ) | ( Ng785  &  (~ n4506) ) ;
 assign Ng24300 = ( (~ n3467) ) ;
 assign n3468 = ( Ng853  &  n343 ) | ( (~ Ng853)  &  (~ Ng488) ) | ( n343  &  (~ Ng488) ) ;
 assign Ng24294 = ( (~ n3468) ) ;
 assign n3469 = ( (~ wire1594)  &  (~ Ng487) ) | ( wire1594  &  n343 ) | ( (~ Ng487)  &  n343 ) ;
 assign Ng24293 = ( (~ n3469) ) ;
 assign n3470 = ( wire1612  &  n343 ) | ( (~ wire1612)  &  (~ Ng486) ) | ( n343  &  (~ Ng486) ) ;
 assign Ng24292 = ( (~ n3470) ) ;
 assign n3471 = ( Ng853  &  (~ n587) ) | ( (~ Ng853)  &  (~ Ng464) ) | ( (~ n587)  &  (~ Ng464) ) ;
 assign Ng24291 = ( (~ n3471) ) ;
 assign n3472 = ( (~ wire1594)  &  (~ Ng484) ) | ( wire1594  &  (~ n587) ) | ( (~ Ng484)  &  (~ n587) ) ;
 assign Ng24290 = ( (~ n3472) ) ;
 assign n3473 = ( wire1612  &  (~ n587) ) | ( (~ wire1612)  &  (~ Ng480) ) | ( (~ n587)  &  (~ Ng480) ) ;
 assign Ng24289 = ( (~ n3473) ) ;
 assign n3474 = ( (~ n613)  &  (~ n2450) ) | ( (~ n613)  &  (~ Ng162) ) | ( n2450  &  (~ Ng162) ) ;
 assign Ng24288 = ( (~ n3474) ) ;
 assign n3475 = ( (~ Ng164)  &  (~ n613) ) | ( (~ Ng164)  &  n4503 ) | ( (~ n613)  &  (~ n4503) ) ;
 assign Ng24287 = ( (~ n3475) ) ;
 assign n3476 = ( (~ n613)  &  (~ Ng163) ) | ( (~ Ng163)  &  n4506 ) | ( (~ n613)  &  (~ n4506) ) ;
 assign Ng24286 = ( (~ n3476) ) ;
 assign n3477 = ( (~ n625)  &  (~ n2450) ) | ( (~ n625)  &  (~ Ng159) ) | ( n2450  &  (~ Ng159) ) ;
 assign Ng24285 = ( (~ n3477) ) ;
 assign n3478 = ( (~ Ng161)  &  (~ n625) ) | ( (~ Ng161)  &  n4503 ) | ( (~ n625)  &  (~ n4503) ) ;
 assign Ng24284 = ( (~ n3478) ) ;
 assign n3479 = ( (~ n625)  &  (~ Ng160) ) | ( (~ Ng160)  &  n4506 ) | ( (~ n625)  &  (~ n4506) ) ;
 assign Ng24283 = ( (~ n3479) ) ;
 assign n3480 = ( Ng125  &  (~ n2450) ) | ( Ng125  &  (~ Ng156) ) | ( n2450  &  (~ Ng156) ) ;
 assign Ng24282 = ( (~ n3480) ) ;
 assign n3481 = ( (~ Ng158)  &  Ng125 ) | ( (~ Ng158)  &  n4503 ) | ( Ng125  &  (~ n4503) ) ;
 assign Ng24281 = ( (~ n3481) ) ;
 assign n3482 = ( Ng125  &  (~ Ng157) ) | ( (~ Ng157)  &  n4506 ) | ( Ng125  &  (~ n4506) ) ;
 assign Ng24280 = ( (~ n3482) ) ;
 assign n3483 = ( Ng121  &  (~ n2450) ) | ( Ng121  &  (~ Ng153) ) | ( n2450  &  (~ Ng153) ) ;
 assign Ng24279 = ( (~ n3483) ) ;
 assign n3484 = ( (~ Ng155)  &  Ng121 ) | ( (~ Ng155)  &  n4503 ) | ( Ng121  &  (~ n4503) ) ;
 assign Ng24278 = ( (~ n3484) ) ;
 assign n3485 = ( Ng121  &  (~ Ng154) ) | ( (~ Ng154)  &  n4506 ) | ( Ng121  &  (~ n4506) ) ;
 assign Ng24277 = ( (~ n3485) ) ;
 assign n3486 = ( Ng117  &  (~ n2450) ) | ( Ng117  &  (~ Ng150) ) | ( n2450  &  (~ Ng150) ) ;
 assign Ng24276 = ( (~ n3486) ) ;
 assign n3487 = ( Ng117  &  (~ Ng152) ) | ( (~ Ng152)  &  n4503 ) | ( Ng117  &  (~ n4503) ) ;
 assign Ng24275 = ( (~ n3487) ) ;
 assign n3488 = ( (~ Ng151)  &  Ng117 ) | ( (~ Ng151)  &  n4506 ) | ( Ng117  &  (~ n4506) ) ;
 assign Ng24274 = ( (~ n3488) ) ;
 assign n3489 = ( Ng113  &  (~ n2450) ) | ( Ng113  &  (~ Ng147) ) | ( n2450  &  (~ Ng147) ) ;
 assign Ng24273 = ( (~ n3489) ) ;
 assign n3490 = ( Ng113  &  (~ Ng149) ) | ( (~ Ng149)  &  n4503 ) | ( Ng113  &  (~ n4503) ) ;
 assign Ng24272 = ( (~ n3490) ) ;
 assign n3491 = ( (~ Ng148)  &  Ng113 ) | ( (~ Ng148)  &  n4506 ) | ( Ng113  &  (~ n4506) ) ;
 assign Ng24271 = ( (~ n3491) ) ;
 assign n3492 = ( Ng109  &  (~ n2450) ) | ( Ng109  &  (~ Ng144) ) | ( n2450  &  (~ Ng144) ) ;
 assign Ng24270 = ( (~ n3492) ) ;
 assign n3493 = ( Ng109  &  (~ Ng146) ) | ( (~ Ng146)  &  n4503 ) | ( Ng109  &  (~ n4503) ) ;
 assign Ng24269 = ( (~ n3493) ) ;
 assign n3494 = ( (~ Ng145)  &  Ng109 ) | ( (~ Ng145)  &  n4506 ) | ( Ng109  &  (~ n4506) ) ;
 assign Ng24268 = ( (~ n3494) ) ;
 assign n3495 = ( Ng105  &  (~ n2450) ) | ( Ng105  &  (~ Ng141) ) | ( n2450  &  (~ Ng141) ) ;
 assign Ng24267 = ( (~ n3495) ) ;
 assign n3496 = ( Ng105  &  (~ Ng143) ) | ( (~ Ng143)  &  n4503 ) | ( Ng105  &  (~ n4503) ) ;
 assign Ng24266 = ( (~ n3496) ) ;
 assign n3497 = ( (~ Ng142)  &  Ng105 ) | ( (~ Ng142)  &  n4506 ) | ( Ng105  &  (~ n4506) ) ;
 assign Ng24265 = ( (~ n3497) ) ;
 assign n3498 = ( Ng101  &  (~ n2450) ) | ( Ng101  &  (~ Ng132) ) | ( n2450  &  (~ Ng132) ) ;
 assign Ng24264 = ( (~ n3498) ) ;
 assign n3499 = ( (~ Ng134)  &  Ng101 ) | ( (~ Ng134)  &  n4503 ) | ( Ng101  &  (~ n4503) ) ;
 assign Ng24263 = ( (~ n3499) ) ;
 assign n3500 = ( Ng101  &  (~ Ng133) ) | ( (~ Ng133)  &  n4506 ) | ( Ng101  &  (~ n4506) ) ;
 assign Ng24262 = ( (~ n3500) ) ;
 assign n3501 = ( Ng97  &  (~ n2450) ) | ( Ng97  &  (~ Ng129) ) | ( n2450  &  (~ Ng129) ) ;
 assign Ng24261 = ( (~ n3501) ) ;
 assign n3502 = ( (~ Ng131)  &  Ng97 ) | ( (~ Ng131)  &  n4503 ) | ( Ng97  &  (~ n4503) ) ;
 assign Ng24260 = ( (~ n3502) ) ;
 assign n3503 = ( Ng97  &  (~ Ng130) ) | ( (~ Ng130)  &  n4506 ) | ( Ng97  &  (~ n4506) ) ;
 assign Ng24259 = ( (~ n3503) ) ;
 assign n3504 = ( (~ Pg8096)  &  Ng2879 ) | ( (~ Pg8096)  &  n4644 ) | ( (~ Ng2879)  &  n4644 ) ;
 assign Ng23316 = ( (~ n3504) ) ;
 assign n3505 = ( (~ Ng2879)  &  (~ Ng13455) ) | ( Ng2879  &  (~ n4900) ) | ( (~ Ng13455)  &  (~ n4900) ) ;
 assign Ng23314 = ( (~ n3505) ) ;
 assign n3506 = ( Ng2879  &  n4644 ) | ( (~ Ng2879)  &  (~ Ng13439) ) | ( n4644  &  (~ Ng13439) ) ;
 assign Ng23313 = ( (~ n3506) ) ;
 assign n3507 = ( (~ Pg7519)  &  Ng2879 ) | ( (~ Pg7519)  &  (~ n4900) ) | ( (~ Ng2879)  &  (~ n4900) ) ;
 assign Ng23312 = ( (~ n3507) ) ;
 assign n3508 = ( (~ n662)  &  (~ n771) ) | ( (~ n662)  &  (~ Ng2805) ) | ( n771  &  (~ Ng2805) ) ;
 assign Ng23311 = ( (~ n3508) ) ;
 assign n3509 = ( (~ Ng2807)  &  (~ n662) ) | ( (~ Ng2807)  &  n713 ) | ( (~ n662)  &  (~ n713) ) ;
 assign Ng23310 = ( (~ n3509) ) ;
 assign n3510 = ( (~ n662)  &  (~ n762) ) | ( (~ n662)  &  (~ Ng2806) ) | ( n762  &  (~ Ng2806) ) ;
 assign Ng23309 = ( (~ n3510) ) ;
 assign n3511 = ( (~ n569)  &  (~ n771) ) | ( (~ n569)  &  (~ Ng2802) ) | ( n771  &  (~ Ng2802) ) ;
 assign Ng23308 = ( (~ n3511) ) ;
 assign n3512 = ( (~ n569)  &  (~ n713) ) | ( (~ n569)  &  (~ Ng2804) ) | ( n713  &  (~ Ng2804) ) ;
 assign Ng23307 = ( (~ n3512) ) ;
 assign n3513 = ( (~ n569)  &  (~ n762) ) | ( (~ n569)  &  (~ Ng2803) ) | ( n762  &  (~ Ng2803) ) ;
 assign Ng23306 = ( (~ n3513) ) ;
 assign n3514 = ( n770  &  Ng2766 ) | ( (~ n770)  &  (~ Ng2799) ) | ( Ng2766  &  (~ Ng2799) ) ;
 assign Ng23305 = ( (~ n3514) ) ;
 assign n3515 = ( (~ Ng2801)  &  (~ n767) ) | ( (~ Ng2801)  &  Ng2766 ) | ( n767  &  Ng2766 ) ;
 assign Ng23304 = ( (~ n3515) ) ;
 assign n3516 = ( n761  &  Ng2766 ) | ( (~ n761)  &  (~ Ng2800) ) | ( Ng2766  &  (~ Ng2800) ) ;
 assign Ng23303 = ( (~ n3516) ) ;
 assign n3517 = ( n770  &  Ng2760 ) | ( (~ n770)  &  (~ Ng2796) ) | ( Ng2760  &  (~ Ng2796) ) ;
 assign Ng23302 = ( (~ n3517) ) ;
 assign n3518 = ( (~ Ng2798)  &  (~ n767) ) | ( (~ Ng2798)  &  Ng2760 ) | ( n767  &  Ng2760 ) ;
 assign Ng23301 = ( (~ n3518) ) ;
 assign n3519 = ( n761  &  Ng2760 ) | ( (~ n761)  &  (~ Ng2797) ) | ( Ng2760  &  (~ Ng2797) ) ;
 assign Ng23300 = ( (~ n3519) ) ;
 assign n3520 = ( n770  &  Ng2753 ) | ( (~ n770)  &  (~ Ng2793) ) | ( Ng2753  &  (~ Ng2793) ) ;
 assign Ng23299 = ( (~ n3520) ) ;
 assign n3521 = ( (~ Ng2795)  &  (~ n767) ) | ( (~ Ng2795)  &  Ng2753 ) | ( n767  &  Ng2753 ) ;
 assign Ng23298 = ( (~ n3521) ) ;
 assign n3522 = ( n761  &  Ng2753 ) | ( (~ n761)  &  (~ Ng2794) ) | ( Ng2753  &  (~ Ng2794) ) ;
 assign Ng23297 = ( (~ n3522) ) ;
 assign n3523 = ( n770  &  Ng2740 ) | ( (~ n770)  &  (~ Ng2790) ) | ( Ng2740  &  (~ Ng2790) ) ;
 assign Ng23296 = ( (~ n3523) ) ;
 assign n3524 = ( (~ Ng2792)  &  (~ n767) ) | ( (~ Ng2792)  &  Ng2740 ) | ( n767  &  Ng2740 ) ;
 assign Ng23295 = ( (~ n3524) ) ;
 assign n3525 = ( n761  &  Ng2740 ) | ( (~ n761)  &  (~ Ng2791) ) | ( Ng2740  &  (~ Ng2791) ) ;
 assign Ng23294 = ( (~ n3525) ) ;
 assign n3526 = ( n770  &  Ng2746 ) | ( (~ n770)  &  (~ Ng2787) ) | ( Ng2746  &  (~ Ng2787) ) ;
 assign Ng23293 = ( (~ n3526) ) ;
 assign n3527 = ( (~ Ng2789)  &  (~ n767) ) | ( (~ Ng2789)  &  Ng2746 ) | ( n767  &  Ng2746 ) ;
 assign Ng23292 = ( (~ n3527) ) ;
 assign n3528 = ( n761  &  Ng2746 ) | ( (~ n761)  &  (~ Ng2788) ) | ( Ng2746  &  (~ Ng2788) ) ;
 assign Ng23291 = ( (~ n3528) ) ;
 assign n3529 = ( n770  &  Ng2734 ) | ( (~ n770)  &  (~ Ng2784) ) | ( Ng2734  &  (~ Ng2784) ) ;
 assign Ng23290 = ( (~ n3529) ) ;
 assign n3530 = ( (~ Ng2786)  &  (~ n767) ) | ( (~ Ng2786)  &  Ng2734 ) | ( n767  &  Ng2734 ) ;
 assign Ng23289 = ( (~ n3530) ) ;
 assign n3531 = ( n761  &  Ng2734 ) | ( (~ n761)  &  (~ Ng2785) ) | ( Ng2734  &  (~ Ng2785) ) ;
 assign Ng23288 = ( (~ n3531) ) ;
 assign n3532 = ( n770  &  Ng2720 ) | ( (~ n770)  &  (~ Ng2781) ) | ( Ng2720  &  (~ Ng2781) ) ;
 assign Ng23287 = ( (~ n3532) ) ;
 assign n3533 = ( (~ Ng2783)  &  (~ n767) ) | ( (~ Ng2783)  &  Ng2720 ) | ( n767  &  Ng2720 ) ;
 assign Ng23286 = ( (~ n3533) ) ;
 assign n3534 = ( n761  &  Ng2720 ) | ( (~ n761)  &  (~ Ng2782) ) | ( Ng2720  &  (~ Ng2782) ) ;
 assign Ng23285 = ( (~ n3534) ) ;
 assign n3535 = ( n770  &  Ng2727 ) | ( (~ n770)  &  (~ Ng2778) ) | ( Ng2727  &  (~ Ng2778) ) ;
 assign Ng23284 = ( (~ n3535) ) ;
 assign n3536 = ( (~ Ng2780)  &  (~ n767) ) | ( (~ Ng2780)  &  Ng2727 ) | ( n767  &  Ng2727 ) ;
 assign Ng23283 = ( (~ n3536) ) ;
 assign n3537 = ( n761  &  Ng2727 ) | ( (~ n761)  &  (~ Ng2779) ) | ( Ng2727  &  (~ Ng2779) ) ;
 assign Ng23282 = ( (~ n3537) ) ;
 assign n3538 = ( n770  &  Ng2707 ) | ( (~ n770)  &  (~ Ng2775) ) | ( Ng2707  &  (~ Ng2775) ) ;
 assign Ng23281 = ( (~ n3538) ) ;
 assign n3539 = ( (~ Ng2777)  &  (~ n767) ) | ( (~ Ng2777)  &  Ng2707 ) | ( n767  &  Ng2707 ) ;
 assign Ng23280 = ( (~ n3539) ) ;
 assign n3540 = ( n761  &  Ng2707 ) | ( (~ n761)  &  (~ Ng2776) ) | ( Ng2707  &  (~ Ng2776) ) ;
 assign Ng23279 = ( (~ n3540) ) ;
 assign n3541 = ( n770  &  Ng2714 ) | ( (~ n770)  &  (~ Ng2772) ) | ( Ng2714  &  (~ Ng2772) ) ;
 assign Ng23278 = ( (~ n3541) ) ;
 assign n3542 = ( (~ Ng2774)  &  (~ n767) ) | ( (~ Ng2774)  &  Ng2714 ) | ( n767  &  Ng2714 ) ;
 assign Ng23277 = ( (~ n3542) ) ;
 assign n3543 = ( n761  &  Ng2714 ) | ( (~ n761)  &  (~ Ng2773) ) | ( Ng2714  &  (~ Ng2773) ) ;
 assign Ng23276 = ( (~ n3543) ) ;
 assign n3544 = ( (~ n659)  &  (~ n766) ) | ( (~ n659)  &  (~ Ng2111) ) | ( n766  &  (~ Ng2111) ) ;
 assign Ng23273 = ( (~ n3544) ) ;
 assign n3545 = ( (~ Ng2113)  &  (~ n659) ) | ( (~ Ng2113)  &  n711 ) | ( (~ n659)  &  (~ n711) ) ;
 assign Ng23272 = ( (~ n3545) ) ;
 assign n3546 = ( (~ n659)  &  (~ n755) ) | ( (~ n659)  &  (~ Ng2112) ) | ( n755  &  (~ Ng2112) ) ;
 assign Ng23271 = ( (~ n3546) ) ;
 assign n3547 = ( (~ n564)  &  (~ n766) ) | ( (~ n564)  &  (~ Ng2108) ) | ( n766  &  (~ Ng2108) ) ;
 assign Ng23270 = ( (~ n3547) ) ;
 assign n3548 = ( (~ n564)  &  (~ n711) ) | ( (~ n564)  &  (~ Ng2110) ) | ( n711  &  (~ Ng2110) ) ;
 assign Ng23269 = ( (~ n3548) ) ;
 assign n3549 = ( (~ n564)  &  (~ n755) ) | ( (~ n564)  &  (~ Ng2109) ) | ( n755  &  (~ Ng2109) ) ;
 assign Ng23268 = ( (~ n3549) ) ;
 assign n3550 = ( n765  &  Ng2072 ) | ( (~ n765)  &  (~ Ng2105) ) | ( Ng2072  &  (~ Ng2105) ) ;
 assign Ng23267 = ( (~ n3550) ) ;
 assign n3551 = ( (~ Ng2107)  &  (~ n760) ) | ( (~ Ng2107)  &  Ng2072 ) | ( n760  &  Ng2072 ) ;
 assign Ng23266 = ( (~ n3551) ) ;
 assign n3552 = ( n754  &  Ng2072 ) | ( (~ n754)  &  (~ Ng2106) ) | ( Ng2072  &  (~ Ng2106) ) ;
 assign Ng23265 = ( (~ n3552) ) ;
 assign n3553 = ( n765  &  Ng2066 ) | ( (~ n765)  &  (~ Ng2102) ) | ( Ng2066  &  (~ Ng2102) ) ;
 assign Ng23264 = ( (~ n3553) ) ;
 assign n3554 = ( (~ Ng2104)  &  (~ n760) ) | ( (~ Ng2104)  &  Ng2066 ) | ( n760  &  Ng2066 ) ;
 assign Ng23263 = ( (~ n3554) ) ;
 assign n3555 = ( n754  &  Ng2066 ) | ( (~ n754)  &  (~ Ng2103) ) | ( Ng2066  &  (~ Ng2103) ) ;
 assign Ng23262 = ( (~ n3555) ) ;
 assign n3556 = ( n765  &  Ng2059 ) | ( (~ n765)  &  (~ Ng2099) ) | ( Ng2059  &  (~ Ng2099) ) ;
 assign Ng23261 = ( (~ n3556) ) ;
 assign n3557 = ( (~ Ng2101)  &  (~ n760) ) | ( (~ Ng2101)  &  Ng2059 ) | ( n760  &  Ng2059 ) ;
 assign Ng23260 = ( (~ n3557) ) ;
 assign n3558 = ( n754  &  Ng2059 ) | ( (~ n754)  &  (~ Ng2100) ) | ( Ng2059  &  (~ Ng2100) ) ;
 assign Ng23259 = ( (~ n3558) ) ;
 assign n3559 = ( n765  &  Ng2046 ) | ( (~ n765)  &  (~ Ng2096) ) | ( Ng2046  &  (~ Ng2096) ) ;
 assign Ng23258 = ( (~ n3559) ) ;
 assign n3560 = ( (~ Ng2098)  &  (~ n760) ) | ( (~ Ng2098)  &  Ng2046 ) | ( n760  &  Ng2046 ) ;
 assign Ng23257 = ( (~ n3560) ) ;
 assign n3561 = ( n754  &  Ng2046 ) | ( (~ n754)  &  (~ Ng2097) ) | ( Ng2046  &  (~ Ng2097) ) ;
 assign Ng23256 = ( (~ n3561) ) ;
 assign n3562 = ( n765  &  Ng2052 ) | ( (~ n765)  &  (~ Ng2093) ) | ( Ng2052  &  (~ Ng2093) ) ;
 assign Ng23255 = ( (~ n3562) ) ;
 assign n3563 = ( (~ Ng2095)  &  (~ n760) ) | ( (~ Ng2095)  &  Ng2052 ) | ( n760  &  Ng2052 ) ;
 assign Ng23254 = ( (~ n3563) ) ;
 assign n3564 = ( n754  &  Ng2052 ) | ( (~ n754)  &  (~ Ng2094) ) | ( Ng2052  &  (~ Ng2094) ) ;
 assign Ng23253 = ( (~ n3564) ) ;
 assign n3565 = ( n765  &  Ng2040 ) | ( (~ n765)  &  (~ Ng2090) ) | ( Ng2040  &  (~ Ng2090) ) ;
 assign Ng23252 = ( (~ n3565) ) ;
 assign n3566 = ( (~ Ng2092)  &  (~ n760) ) | ( (~ Ng2092)  &  Ng2040 ) | ( n760  &  Ng2040 ) ;
 assign Ng23251 = ( (~ n3566) ) ;
 assign n3567 = ( n754  &  Ng2040 ) | ( (~ n754)  &  (~ Ng2091) ) | ( Ng2040  &  (~ Ng2091) ) ;
 assign Ng23250 = ( (~ n3567) ) ;
 assign n3568 = ( n765  &  Ng2026 ) | ( (~ n765)  &  (~ Ng2087) ) | ( Ng2026  &  (~ Ng2087) ) ;
 assign Ng23249 = ( (~ n3568) ) ;
 assign n3569 = ( (~ Ng2089)  &  (~ n760) ) | ( (~ Ng2089)  &  Ng2026 ) | ( n760  &  Ng2026 ) ;
 assign Ng23248 = ( (~ n3569) ) ;
 assign n3570 = ( n754  &  Ng2026 ) | ( (~ n754)  &  (~ Ng2088) ) | ( Ng2026  &  (~ Ng2088) ) ;
 assign Ng23247 = ( (~ n3570) ) ;
 assign n3571 = ( n765  &  Ng2033 ) | ( (~ n765)  &  (~ Ng2084) ) | ( Ng2033  &  (~ Ng2084) ) ;
 assign Ng23246 = ( (~ n3571) ) ;
 assign n3572 = ( (~ Ng2086)  &  (~ n760) ) | ( (~ Ng2086)  &  Ng2033 ) | ( n760  &  Ng2033 ) ;
 assign Ng23245 = ( (~ n3572) ) ;
 assign n3573 = ( n754  &  Ng2033 ) | ( (~ n754)  &  (~ Ng2085) ) | ( Ng2033  &  (~ Ng2085) ) ;
 assign Ng23244 = ( (~ n3573) ) ;
 assign n3574 = ( n765  &  Ng2013 ) | ( (~ n765)  &  (~ Ng2081) ) | ( Ng2013  &  (~ Ng2081) ) ;
 assign Ng23243 = ( (~ n3574) ) ;
 assign n3575 = ( (~ Ng2083)  &  (~ n760) ) | ( (~ Ng2083)  &  Ng2013 ) | ( n760  &  Ng2013 ) ;
 assign Ng23242 = ( (~ n3575) ) ;
 assign n3576 = ( n754  &  Ng2013 ) | ( (~ n754)  &  (~ Ng2082) ) | ( Ng2013  &  (~ Ng2082) ) ;
 assign Ng23241 = ( (~ n3576) ) ;
 assign n3577 = ( n765  &  Ng2020 ) | ( (~ n765)  &  (~ Ng2078) ) | ( Ng2020  &  (~ Ng2078) ) ;
 assign Ng23240 = ( (~ n3577) ) ;
 assign n3578 = ( (~ Ng2080)  &  (~ n760) ) | ( (~ Ng2080)  &  Ng2020 ) | ( n760  &  Ng2020 ) ;
 assign Ng23239 = ( (~ n3578) ) ;
 assign n3579 = ( n754  &  Ng2020 ) | ( (~ n754)  &  (~ Ng2079) ) | ( Ng2020  &  (~ Ng2079) ) ;
 assign Ng23238 = ( (~ n3579) ) ;
 assign n3580 = ( (~ n654)  &  (~ n759) ) | ( (~ n654)  &  (~ Ng1417) ) | ( n759  &  (~ Ng1417) ) ;
 assign Ng23235 = ( (~ n3580) ) ;
 assign n3581 = ( (~ Ng1419)  &  (~ n654) ) | ( (~ Ng1419)  &  n709 ) | ( (~ n654)  &  (~ n709) ) ;
 assign Ng23234 = ( (~ n3581) ) ;
 assign n3582 = ( (~ n654)  &  (~ n748) ) | ( (~ n654)  &  (~ Ng1418) ) | ( n748  &  (~ Ng1418) ) ;
 assign Ng23233 = ( (~ n3582) ) ;
 assign n3583 = ( (~ n557)  &  (~ n759) ) | ( (~ n557)  &  (~ Ng1414) ) | ( n759  &  (~ Ng1414) ) ;
 assign Ng23232 = ( (~ n3583) ) ;
 assign n3584 = ( (~ n557)  &  (~ n709) ) | ( (~ n557)  &  (~ Ng1416) ) | ( n709  &  (~ Ng1416) ) ;
 assign Ng23231 = ( (~ n3584) ) ;
 assign n3585 = ( (~ n557)  &  (~ n748) ) | ( (~ n557)  &  (~ Ng1415) ) | ( n748  &  (~ Ng1415) ) ;
 assign Ng23230 = ( (~ n3585) ) ;
 assign n3586 = ( n758  &  Ng1378 ) | ( (~ n758)  &  (~ Ng1411) ) | ( Ng1378  &  (~ Ng1411) ) ;
 assign Ng23229 = ( (~ n3586) ) ;
 assign n3587 = ( (~ Ng1413)  &  (~ n753) ) | ( (~ Ng1413)  &  Ng1378 ) | ( n753  &  Ng1378 ) ;
 assign Ng23228 = ( (~ n3587) ) ;
 assign n3588 = ( n747  &  Ng1378 ) | ( (~ n747)  &  (~ Ng1412) ) | ( Ng1378  &  (~ Ng1412) ) ;
 assign Ng23227 = ( (~ n3588) ) ;
 assign n3589 = ( n758  &  Ng1372 ) | ( (~ n758)  &  (~ Ng1408) ) | ( Ng1372  &  (~ Ng1408) ) ;
 assign Ng23226 = ( (~ n3589) ) ;
 assign n3590 = ( (~ Ng1410)  &  (~ n753) ) | ( (~ Ng1410)  &  Ng1372 ) | ( n753  &  Ng1372 ) ;
 assign Ng23225 = ( (~ n3590) ) ;
 assign n3591 = ( n747  &  Ng1372 ) | ( (~ n747)  &  (~ Ng1409) ) | ( Ng1372  &  (~ Ng1409) ) ;
 assign Ng23224 = ( (~ n3591) ) ;
 assign n3592 = ( n758  &  Ng1365 ) | ( (~ n758)  &  (~ Ng1405) ) | ( Ng1365  &  (~ Ng1405) ) ;
 assign Ng23223 = ( (~ n3592) ) ;
 assign n3593 = ( (~ Ng1407)  &  (~ n753) ) | ( (~ Ng1407)  &  Ng1365 ) | ( n753  &  Ng1365 ) ;
 assign Ng23222 = ( (~ n3593) ) ;
 assign n3594 = ( n747  &  Ng1365 ) | ( (~ n747)  &  (~ Ng1406) ) | ( Ng1365  &  (~ Ng1406) ) ;
 assign Ng23221 = ( (~ n3594) ) ;
 assign n3595 = ( n758  &  Ng1352 ) | ( (~ n758)  &  (~ Ng1402) ) | ( Ng1352  &  (~ Ng1402) ) ;
 assign Ng23220 = ( (~ n3595) ) ;
 assign n3596 = ( (~ Ng1404)  &  (~ n753) ) | ( (~ Ng1404)  &  Ng1352 ) | ( n753  &  Ng1352 ) ;
 assign Ng23219 = ( (~ n3596) ) ;
 assign n3597 = ( n747  &  Ng1352 ) | ( (~ n747)  &  (~ Ng1403) ) | ( Ng1352  &  (~ Ng1403) ) ;
 assign Ng23218 = ( (~ n3597) ) ;
 assign n3598 = ( n758  &  Ng1358 ) | ( (~ n758)  &  (~ Ng1399) ) | ( Ng1358  &  (~ Ng1399) ) ;
 assign Ng23217 = ( (~ n3598) ) ;
 assign n3599 = ( (~ Ng1401)  &  (~ n753) ) | ( (~ Ng1401)  &  Ng1358 ) | ( n753  &  Ng1358 ) ;
 assign Ng23216 = ( (~ n3599) ) ;
 assign n3600 = ( n747  &  Ng1358 ) | ( (~ n747)  &  (~ Ng1400) ) | ( Ng1358  &  (~ Ng1400) ) ;
 assign Ng23215 = ( (~ n3600) ) ;
 assign n3601 = ( n758  &  Ng1346 ) | ( (~ n758)  &  (~ Ng1396) ) | ( Ng1346  &  (~ Ng1396) ) ;
 assign Ng23214 = ( (~ n3601) ) ;
 assign n3602 = ( (~ Ng1398)  &  (~ n753) ) | ( (~ Ng1398)  &  Ng1346 ) | ( n753  &  Ng1346 ) ;
 assign Ng23213 = ( (~ n3602) ) ;
 assign n3603 = ( n747  &  Ng1346 ) | ( (~ n747)  &  (~ Ng1397) ) | ( Ng1346  &  (~ Ng1397) ) ;
 assign Ng23212 = ( (~ n3603) ) ;
 assign n3604 = ( n758  &  Ng1332 ) | ( (~ n758)  &  (~ Ng1393) ) | ( Ng1332  &  (~ Ng1393) ) ;
 assign Ng23211 = ( (~ n3604) ) ;
 assign n3605 = ( (~ Ng1395)  &  (~ n753) ) | ( (~ Ng1395)  &  Ng1332 ) | ( n753  &  Ng1332 ) ;
 assign Ng23210 = ( (~ n3605) ) ;
 assign n3606 = ( n747  &  Ng1332 ) | ( (~ n747)  &  (~ Ng1394) ) | ( Ng1332  &  (~ Ng1394) ) ;
 assign Ng23209 = ( (~ n3606) ) ;
 assign n3607 = ( n758  &  Ng1339 ) | ( (~ n758)  &  (~ Ng1390) ) | ( Ng1339  &  (~ Ng1390) ) ;
 assign Ng23208 = ( (~ n3607) ) ;
 assign n3608 = ( (~ Ng1392)  &  (~ n753) ) | ( (~ Ng1392)  &  Ng1339 ) | ( n753  &  Ng1339 ) ;
 assign Ng23207 = ( (~ n3608) ) ;
 assign n3609 = ( n747  &  Ng1339 ) | ( (~ n747)  &  (~ Ng1391) ) | ( Ng1339  &  (~ Ng1391) ) ;
 assign Ng23206 = ( (~ n3609) ) ;
 assign n3610 = ( n758  &  Ng1319 ) | ( (~ n758)  &  (~ Ng1387) ) | ( Ng1319  &  (~ Ng1387) ) ;
 assign Ng23205 = ( (~ n3610) ) ;
 assign n3611 = ( (~ Ng1389)  &  (~ n753) ) | ( (~ Ng1389)  &  Ng1319 ) | ( n753  &  Ng1319 ) ;
 assign Ng23204 = ( (~ n3611) ) ;
 assign n3612 = ( n747  &  Ng1319 ) | ( (~ n747)  &  (~ Ng1388) ) | ( Ng1319  &  (~ Ng1388) ) ;
 assign Ng23203 = ( (~ n3612) ) ;
 assign n3613 = ( n758  &  Ng1326 ) | ( (~ n758)  &  (~ Ng1384) ) | ( Ng1326  &  (~ Ng1384) ) ;
 assign Ng23202 = ( (~ n3613) ) ;
 assign n3614 = ( (~ Ng1386)  &  (~ n753) ) | ( (~ Ng1386)  &  Ng1326 ) | ( n753  &  Ng1326 ) ;
 assign Ng23201 = ( (~ n3614) ) ;
 assign n3615 = ( n747  &  Ng1326 ) | ( (~ n747)  &  (~ Ng1385) ) | ( Ng1326  &  (~ Ng1385) ) ;
 assign Ng23200 = ( (~ n3615) ) ;
 assign n3616 = ( (~ n649)  &  (~ n752) ) | ( (~ n649)  &  (~ Ng731) ) | ( n752  &  (~ Ng731) ) ;
 assign Ng23197 = ( (~ n3616) ) ;
 assign n3617 = ( (~ Ng733)  &  (~ n649) ) | ( (~ Ng733)  &  n707 ) | ( (~ n649)  &  (~ n707) ) ;
 assign Ng23196 = ( (~ n3617) ) ;
 assign n3618 = ( (~ n649)  &  (~ n744) ) | ( (~ n649)  &  (~ Ng732) ) | ( n744  &  (~ Ng732) ) ;
 assign Ng23195 = ( (~ n3618) ) ;
 assign n3619 = ( (~ n548)  &  (~ n752) ) | ( (~ n548)  &  (~ Ng728) ) | ( n752  &  (~ Ng728) ) ;
 assign Ng23194 = ( (~ n3619) ) ;
 assign n3620 = ( (~ n548)  &  (~ n707) ) | ( (~ n548)  &  (~ Ng730) ) | ( n707  &  (~ Ng730) ) ;
 assign Ng23193 = ( (~ n3620) ) ;
 assign n3621 = ( (~ n548)  &  (~ n744) ) | ( (~ n548)  &  (~ Ng729) ) | ( n744  &  (~ Ng729) ) ;
 assign Ng23192 = ( (~ n3621) ) ;
 assign n3622 = ( n751  &  Ng692 ) | ( (~ n751)  &  (~ Ng725) ) | ( Ng692  &  (~ Ng725) ) ;
 assign Ng23191 = ( (~ n3622) ) ;
 assign n3623 = ( (~ Ng727)  &  (~ n746) ) | ( (~ Ng727)  &  Ng692 ) | ( n746  &  Ng692 ) ;
 assign Ng23190 = ( (~ n3623) ) ;
 assign n3624 = ( n743  &  Ng692 ) | ( (~ n743)  &  (~ Ng726) ) | ( Ng692  &  (~ Ng726) ) ;
 assign Ng23189 = ( (~ n3624) ) ;
 assign n3625 = ( n751  &  Ng686 ) | ( (~ n751)  &  (~ Ng722) ) | ( Ng686  &  (~ Ng722) ) ;
 assign Ng23188 = ( (~ n3625) ) ;
 assign n3626 = ( (~ Ng724)  &  (~ n746) ) | ( (~ Ng724)  &  Ng686 ) | ( n746  &  Ng686 ) ;
 assign Ng23187 = ( (~ n3626) ) ;
 assign n3627 = ( n743  &  Ng686 ) | ( (~ n743)  &  (~ Ng723) ) | ( Ng686  &  (~ Ng723) ) ;
 assign Ng23186 = ( (~ n3627) ) ;
 assign n3628 = ( n751  &  Ng679 ) | ( (~ n751)  &  (~ Ng719) ) | ( Ng679  &  (~ Ng719) ) ;
 assign Ng23185 = ( (~ n3628) ) ;
 assign n3629 = ( (~ Ng721)  &  (~ n746) ) | ( (~ Ng721)  &  Ng679 ) | ( n746  &  Ng679 ) ;
 assign Ng23184 = ( (~ n3629) ) ;
 assign n3630 = ( n743  &  Ng679 ) | ( (~ n743)  &  (~ Ng720) ) | ( Ng679  &  (~ Ng720) ) ;
 assign Ng23183 = ( (~ n3630) ) ;
 assign n3631 = ( n751  &  Ng666 ) | ( (~ n751)  &  (~ Ng716) ) | ( Ng666  &  (~ Ng716) ) ;
 assign Ng23182 = ( (~ n3631) ) ;
 assign n3632 = ( (~ Ng718)  &  (~ n746) ) | ( (~ Ng718)  &  Ng666 ) | ( n746  &  Ng666 ) ;
 assign Ng23181 = ( (~ n3632) ) ;
 assign n3633 = ( n743  &  Ng666 ) | ( (~ n743)  &  (~ Ng717) ) | ( Ng666  &  (~ Ng717) ) ;
 assign Ng23180 = ( (~ n3633) ) ;
 assign n3634 = ( n751  &  Ng672 ) | ( (~ n751)  &  (~ Ng713) ) | ( Ng672  &  (~ Ng713) ) ;
 assign Ng23179 = ( (~ n3634) ) ;
 assign n3635 = ( (~ Ng715)  &  (~ n746) ) | ( (~ Ng715)  &  Ng672 ) | ( n746  &  Ng672 ) ;
 assign Ng23178 = ( (~ n3635) ) ;
 assign n3636 = ( n743  &  Ng672 ) | ( (~ n743)  &  (~ Ng714) ) | ( Ng672  &  (~ Ng714) ) ;
 assign Ng23177 = ( (~ n3636) ) ;
 assign n3637 = ( n751  &  Ng660 ) | ( (~ n751)  &  (~ Ng710) ) | ( Ng660  &  (~ Ng710) ) ;
 assign Ng23176 = ( (~ n3637) ) ;
 assign n3638 = ( (~ Ng712)  &  (~ n746) ) | ( (~ Ng712)  &  Ng660 ) | ( n746  &  Ng660 ) ;
 assign Ng23175 = ( (~ n3638) ) ;
 assign n3639 = ( n743  &  Ng660 ) | ( (~ n743)  &  (~ Ng711) ) | ( Ng660  &  (~ Ng711) ) ;
 assign Ng23174 = ( (~ n3639) ) ;
 assign n3640 = ( n751  &  Ng646 ) | ( (~ n751)  &  (~ Ng707) ) | ( Ng646  &  (~ Ng707) ) ;
 assign Ng23173 = ( (~ n3640) ) ;
 assign n3641 = ( (~ Ng709)  &  (~ n746) ) | ( (~ Ng709)  &  Ng646 ) | ( n746  &  Ng646 ) ;
 assign Ng23172 = ( (~ n3641) ) ;
 assign n3642 = ( n743  &  Ng646 ) | ( (~ n743)  &  (~ Ng708) ) | ( Ng646  &  (~ Ng708) ) ;
 assign Ng23171 = ( (~ n3642) ) ;
 assign n3643 = ( n751  &  Ng653 ) | ( (~ n751)  &  (~ Ng704) ) | ( Ng653  &  (~ Ng704) ) ;
 assign Ng23170 = ( (~ n3643) ) ;
 assign n3644 = ( (~ Ng706)  &  (~ n746) ) | ( (~ Ng706)  &  Ng653 ) | ( n746  &  Ng653 ) ;
 assign Ng23169 = ( (~ n3644) ) ;
 assign n3645 = ( n743  &  Ng653 ) | ( (~ n743)  &  (~ Ng705) ) | ( Ng653  &  (~ Ng705) ) ;
 assign Ng23168 = ( (~ n3645) ) ;
 assign n3646 = ( n751  &  Ng633 ) | ( (~ n751)  &  (~ Ng701) ) | ( Ng633  &  (~ Ng701) ) ;
 assign Ng23167 = ( (~ n3646) ) ;
 assign n3647 = ( (~ Ng703)  &  (~ n746) ) | ( (~ Ng703)  &  Ng633 ) | ( n746  &  Ng633 ) ;
 assign Ng23166 = ( (~ n3647) ) ;
 assign n3648 = ( n743  &  Ng633 ) | ( (~ n743)  &  (~ Ng702) ) | ( Ng633  &  (~ Ng702) ) ;
 assign Ng23165 = ( (~ n3648) ) ;
 assign n3649 = ( n751  &  Ng640 ) | ( (~ n751)  &  (~ Ng698) ) | ( Ng640  &  (~ Ng698) ) ;
 assign Ng23164 = ( (~ n3649) ) ;
 assign n3650 = ( (~ Ng700)  &  (~ n746) ) | ( (~ Ng700)  &  Ng640 ) | ( n746  &  Ng640 ) ;
 assign Ng23163 = ( (~ n3650) ) ;
 assign n3651 = ( n743  &  Ng640 ) | ( (~ n743)  &  (~ Ng699) ) | ( Ng640  &  (~ Ng699) ) ;
 assign Ng23162 = ( (~ n3651) ) ;
 assign n3652 = ( (~ Pg4590)  &  Ng2879 ) | ( (~ Pg4590)  &  (~ Ng2975) ) | ( (~ Ng2879)  &  (~ Ng2975) ) ;
 assign Ng21963 = ( (~ n3652) ) ;
 assign n3653 = ( (~ Pg4323)  &  Ng2879 ) | ( (~ Pg4323)  &  (~ Ng2978) ) | ( (~ Ng2879)  &  (~ Ng2978) ) ;
 assign Ng21962 = ( (~ n3653) ) ;
 assign n3654 = ( (~ Pg4090)  &  Ng2879 ) | ( (~ Pg4090)  &  (~ Ng2981) ) | ( (~ Ng2879)  &  (~ Ng2981) ) ;
 assign Ng21961 = ( (~ n3654) ) ;
 assign n3655 = ( (~ Pg8251)  &  Ng2879 ) | ( (~ Pg8251)  &  (~ Ng2874) ) | ( (~ Ng2879)  &  (~ Ng2874) ) ;
 assign Ng21960 = ( (~ n3655) ) ;
 assign n3656 = ( (~ Pg4450)  &  Ng2879 ) | ( (~ Pg4450)  &  (~ Ng2935) ) | ( (~ Ng2879)  &  (~ Ng2935) ) ;
 assign Ng21959 = ( (~ n3656) ) ;
 assign n3657 = ( (~ Pg4200)  &  Ng2879 ) | ( (~ Pg4200)  &  (~ Ng2938) ) | ( (~ Ng2879)  &  (~ Ng2938) ) ;
 assign Ng21958 = ( (~ n3657) ) ;
 assign n3658 = ( (~ Pg3993)  &  Ng2879 ) | ( (~ Pg3993)  &  (~ Ng2941) ) | ( (~ Ng2879)  &  (~ Ng2941) ) ;
 assign Ng21957 = ( (~ n3658) ) ;
 assign n3659 = ( (~ Pg8175)  &  Ng2879 ) | ( (~ Pg8175)  &  (~ Ng2944) ) | ( (~ Ng2879)  &  (~ Ng2944) ) ;
 assign Ng21956 = ( (~ n3659) ) ;
 assign n3660 = ( (~ Pg8023)  &  Ng2879 ) | ( (~ Pg8023)  &  (~ Ng2947) ) | ( (~ Ng2879)  &  (~ Ng2947) ) ;
 assign Ng21955 = ( (~ n3660) ) ;
 assign n3661 = ( (~ Pg4321)  &  Ng2879 ) | ( (~ Pg4321)  &  (~ Ng2953) ) | ( (~ Ng2879)  &  (~ Ng2953) ) ;
 assign Ng21954 = ( (~ n3661) ) ;
 assign n3662 = ( (~ Pg4088)  &  Ng2879 ) | ( (~ Pg4088)  &  (~ Ng2956) ) | ( (~ Ng2879)  &  (~ Ng2956) ) ;
 assign Ng21953 = ( (~ n3662) ) ;
 assign n3663 = ( (~ Pg8249)  &  Ng2879 ) | ( (~ Pg8249)  &  (~ Ng2959) ) | ( (~ Ng2879)  &  (~ Ng2959) ) ;
 assign Ng21952 = ( (~ n3663) ) ;
 assign n3664 = ( (~ Pg7334)  &  Ng2879 ) | ( (~ Pg7334)  &  (~ Ng2963) ) | ( (~ Ng2879)  &  (~ Ng2963) ) ;
 assign Ng21950 = ( (~ n3664) ) ;
 assign n3665 = ( (~ Pg6895)  &  Ng2879 ) | ( (~ Pg6895)  &  (~ Ng2966) ) | ( (~ Ng2879)  &  (~ Ng2966) ) ;
 assign Ng21949 = ( (~ n3665) ) ;
 assign n3666 = ( (~ Pg6442)  &  Ng2879 ) | ( (~ Pg6442)  &  (~ Ng2969) ) | ( (~ Ng2879)  &  (~ Ng2969) ) ;
 assign Ng21948 = ( (~ n3666) ) ;
 assign n3667 = ( (~ Pg6225)  &  Ng2879 ) | ( (~ Pg6225)  &  (~ Ng2972) ) | ( (~ Ng2879)  &  (~ Ng2972) ) ;
 assign Ng21947 = ( (~ n3667) ) ;
 assign n3668 = ( Ng1315  &  (~ Ng559) ) | ( (~ Ng1315)  &  (~ Ng3084) ) | ( (~ Ng559)  &  (~ Ng3084) ) ;
 assign Ng20632 = ( (~ n3668) ) ;
 assign n3669 = ( wire1603  &  (~ Ng559) ) | ( (~ wire1603)  &  (~ Ng3211) ) | ( (~ Ng559)  &  (~ Ng3211) ) ;
 assign Ng20631 = ( (~ n3669) ) ;
 assign n3670 = ( wire1605  &  (~ Ng559) ) | ( (~ wire1605)  &  (~ Ng3210) ) | ( (~ Ng559)  &  (~ Ng3210) ) ;
 assign Ng20630 = ( (~ n3670) ) ;
 assign n3671 = ( Ng1315  &  (~ Ng8311) ) | ( (~ Ng1315)  &  (~ Ng3088) ) | ( (~ Ng8311)  &  (~ Ng3088) ) ;
 assign Ng20629 = ( (~ n3671) ) ;
 assign n3672 = ( wire1603  &  (~ Ng8311) ) | ( (~ wire1603)  &  (~ Ng3185) ) | ( (~ Ng8311)  &  (~ Ng3185) ) ;
 assign Ng20628 = ( (~ n3672) ) ;
 assign n3673 = ( wire1605  &  (~ Ng8311) ) | ( (~ wire1605)  &  (~ Ng3182) ) | ( (~ Ng8311)  &  (~ Ng3182) ) ;
 assign Ng20627 = ( (~ n3673) ) ;
 assign n3674 = ( Ng1315  &  (~ Ng8302) ) | ( (~ Ng1315)  &  (~ Ng3179) ) | ( (~ Ng8302)  &  (~ Ng3179) ) ;
 assign Ng20626 = ( (~ n3674) ) ;
 assign n3675 = ( wire1603  &  (~ Ng8302) ) | ( (~ wire1603)  &  (~ Ng3176) ) | ( (~ Ng8302)  &  (~ Ng3176) ) ;
 assign Ng20625 = ( (~ n3675) ) ;
 assign n3676 = ( wire1605  &  (~ Ng8302) ) | ( (~ wire1605)  &  (~ Ng3173) ) | ( (~ Ng8302)  &  (~ Ng3173) ) ;
 assign Ng20624 = ( (~ n3676) ) ;
 assign n3677 = ( Ng1315  &  (~ Ng8293) ) | ( (~ Ng1315)  &  (~ Ng3170) ) | ( (~ Ng8293)  &  (~ Ng3170) ) ;
 assign Ng20623 = ( (~ n3677) ) ;
 assign n3678 = ( wire1603  &  (~ Ng8293) ) | ( (~ wire1603)  &  (~ Ng3167) ) | ( (~ Ng8293)  &  (~ Ng3167) ) ;
 assign Ng20622 = ( (~ n3678) ) ;
 assign n3679 = ( wire1605  &  (~ Ng8293) ) | ( (~ wire1605)  &  (~ Ng3164) ) | ( (~ Ng8293)  &  (~ Ng3164) ) ;
 assign Ng20621 = ( (~ n3679) ) ;
 assign n3680 = ( Ng1315  &  (~ Ng8284) ) | ( (~ Ng1315)  &  (~ Ng3161) ) | ( (~ Ng8284)  &  (~ Ng3161) ) ;
 assign Ng20620 = ( (~ n3680) ) ;
 assign n3681 = ( wire1603  &  (~ Ng8284) ) | ( (~ wire1603)  &  (~ Ng3158) ) | ( (~ Ng8284)  &  (~ Ng3158) ) ;
 assign Ng20619 = ( (~ n3681) ) ;
 assign n3682 = ( wire1605  &  (~ Ng8284) ) | ( (~ wire1605)  &  (~ Ng3155) ) | ( (~ Ng8284)  &  (~ Ng3155) ) ;
 assign Ng20618 = ( (~ n3682) ) ;
 assign n3683 = ( Ng1315  &  (~ Ng2633) ) | ( (~ Ng1315)  &  (~ Ng3096) ) | ( (~ Ng2633)  &  (~ Ng3096) ) ;
 assign Ng20617 = ( (~ n3683) ) ;
 assign n3684 = ( wire1603  &  (~ Ng2633) ) | ( (~ wire1603)  &  (~ Ng3095) ) | ( (~ Ng2633)  &  (~ Ng3095) ) ;
 assign Ng20616 = ( (~ n3684) ) ;
 assign n3685 = ( wire1605  &  (~ Ng2633) ) | ( (~ wire1605)  &  (~ Ng3094) ) | ( (~ Ng2633)  &  (~ Ng3094) ) ;
 assign Ng20615 = ( (~ n3685) ) ;
 assign n3686 = ( Ng1315  &  (~ Ng1939) ) | ( (~ Ng1315)  &  (~ Ng3093) ) | ( (~ Ng1939)  &  (~ Ng3093) ) ;
 assign Ng20614 = ( (~ n3686) ) ;
 assign n3687 = ( wire1603  &  (~ Ng1939) ) | ( (~ wire1603)  &  (~ Ng3092) ) | ( (~ Ng1939)  &  (~ Ng3092) ) ;
 assign Ng20613 = ( (~ n3687) ) ;
 assign n3688 = ( wire1605  &  (~ Ng1939) ) | ( (~ wire1605)  &  (~ Ng3091) ) | ( (~ Ng1939)  &  (~ Ng3091) ) ;
 assign Ng20612 = ( (~ n3688) ) ;
 assign n3689 = ( Ng1315  &  (~ Ng1245) ) | ( (~ Ng1315)  &  (~ Ng3087) ) | ( (~ Ng1245)  &  (~ Ng3087) ) ;
 assign Ng20611 = ( (~ n3689) ) ;
 assign n3690 = ( wire1603  &  (~ Ng1245) ) | ( (~ wire1603)  &  (~ Ng3086) ) | ( (~ Ng1245)  &  (~ Ng3086) ) ;
 assign Ng20610 = ( (~ n3690) ) ;
 assign n3691 = ( wire1605  &  (~ Ng1245) ) | ( (~ wire1605)  &  (~ Ng3085) ) | ( (~ Ng1245)  &  (~ Ng3085) ) ;
 assign Ng20609 = ( (~ n3691) ) ;
 assign n3692 = ( (~ Ng2987)  &  (~ Ng3056) ) | ( Ng2987  &  (~ Ng3074) ) | ( (~ Ng3056)  &  (~ Ng3074) ) ;
 assign Ng20608 = ( (~ n3692) ) ;
 assign n3693 = ( (~ Ng2987)  &  (~ Ng3055) ) | ( Ng2987  &  (~ Ng3073) ) | ( (~ Ng3055)  &  (~ Ng3073) ) ;
 assign Ng20607 = ( (~ n3693) ) ;
 assign n3694 = ( (~ Ng2987)  &  (~ Ng3053) ) | ( Ng2987  &  (~ Ng3072) ) | ( (~ Ng3053)  &  (~ Ng3072) ) ;
 assign Ng20606 = ( (~ n3694) ) ;
 assign n3695 = ( (~ Ng2987)  &  (~ Ng3052) ) | ( Ng2987  &  (~ Ng3071) ) | ( (~ Ng3052)  &  (~ Ng3071) ) ;
 assign Ng20605 = ( (~ n3695) ) ;
 assign n3696 = ( (~ Ng2987)  &  (~ Ng3051) ) | ( Ng2987  &  (~ Ng3070) ) | ( (~ Ng3051)  &  (~ Ng3070) ) ;
 assign Ng20603 = ( (~ n3696) ) ;
 assign n3697 = ( (~ Ng2987)  &  (~ Ng3050) ) | ( Ng2987  &  (~ Ng3069) ) | ( (~ Ng3050)  &  (~ Ng3069) ) ;
 assign Ng20602 = ( (~ n3697) ) ;
 assign n3698 = ( (~ Ng2987)  &  (~ Ng3049) ) | ( Ng2987  &  (~ Ng3068) ) | ( (~ Ng3049)  &  (~ Ng3068) ) ;
 assign Ng20601 = ( (~ n3698) ) ;
 assign n3699 = ( (~ Ng2987)  &  (~ Ng3048) ) | ( Ng2987  &  (~ Ng3067) ) | ( (~ Ng3048)  &  (~ Ng3067) ) ;
 assign Ng20600 = ( (~ n3699) ) ;
 assign n3700 = ( (~ Ng2987)  &  (~ Ng3047) ) | ( Ng2987  &  (~ Ng3066) ) | ( (~ Ng3047)  &  (~ Ng3066) ) ;
 assign Ng20599 = ( (~ n3700) ) ;
 assign n3701 = ( (~ Ng2987)  &  (~ Ng3046) ) | ( Ng2987  &  (~ Ng3065) ) | ( (~ Ng3046)  &  (~ Ng3065) ) ;
 assign Ng20598 = ( (~ n3701) ) ;
 assign n3702 = ( (~ Ng2987)  &  (~ Ng3045) ) | ( Ng2987  &  (~ Ng3064) ) | ( (~ Ng3045)  &  (~ Ng3064) ) ;
 assign Ng20597 = ( (~ n3702) ) ;
 assign n3703 = ( (~ Ng2987)  &  (~ Ng3044) ) | ( Ng2987  &  (~ Ng3063) ) | ( (~ Ng3044)  &  (~ Ng3063) ) ;
 assign Ng20596 = ( (~ n3703) ) ;
 assign n3704 = ( (~ Ng2987)  &  (~ Ng3043) ) | ( Ng2987  &  (~ Ng3062) ) | ( (~ Ng3043)  &  (~ Ng3062) ) ;
 assign Ng20595 = ( (~ n3704) ) ;
 assign n3705 = ( (~ Ng2987)  &  (~ Ng3061) ) | ( Ng2987  &  (~ Ng2997) ) | ( (~ Ng3061)  &  (~ Ng2997) ) ;
 assign Ng20593 = ( (~ n3705) ) ;
 assign n3706 = ( (~ Ng2987)  &  (~ Ng3060) ) | ( Ng2987  &  (~ Ng3078) ) | ( (~ Ng3060)  &  (~ Ng3078) ) ;
 assign Ng20592 = ( (~ n3706) ) ;
 assign n3707 = ( (~ Ng2987)  &  (~ Ng3059) ) | ( Ng2987  &  (~ Ng3077) ) | ( (~ Ng3059)  &  (~ Ng3077) ) ;
 assign Ng20591 = ( (~ n3707) ) ;
 assign n3708 = ( (~ Ng2987)  &  (~ Ng3058) ) | ( Ng2987  &  (~ Ng3076) ) | ( (~ Ng3058)  &  (~ Ng3076) ) ;
 assign Ng20590 = ( (~ n3708) ) ;
 assign n3709 = ( (~ Ng2987)  &  (~ Ng3057) ) | ( Ng2987  &  (~ Ng3075) ) | ( (~ Ng3057)  &  (~ Ng3075) ) ;
 assign Ng20589 = ( (~ n3709) ) ;
 assign n3710 = ( (~ Ng2200)  &  (~ Ng2879) ) | ( (~ Ng2200)  &  (~ Ng2874) ) | ( Ng2879  &  (~ Ng2874) ) ;
 assign Ng20587 = ( (~ n3710) ) ;
 assign n3711 = ( (~ Ng2190)  &  (~ Ng2879) ) | ( (~ Ng2190)  &  (~ Ng2978) ) | ( Ng2879  &  (~ Ng2978) ) ;
 assign Ng20586 = ( (~ n3711) ) ;
 assign n3712 = ( (~ Ng2195)  &  (~ Ng2879) ) | ( (~ Ng2195)  &  (~ Ng2981) ) | ( Ng2879  &  (~ Ng2981) ) ;
 assign Ng20585 = ( (~ n3712) ) ;
 assign n3713 = ( (~ Ng2185)  &  (~ Ng2879) ) | ( (~ Ng2185)  &  (~ Ng2975) ) | ( Ng2879  &  (~ Ng2975) ) ;
 assign Ng20584 = ( (~ n3713) ) ;
 assign n3714 = ( (~ Ng2180)  &  (~ Ng2879) ) | ( (~ Ng2180)  &  (~ Ng2972) ) | ( Ng2879  &  (~ Ng2972) ) ;
 assign Ng20583 = ( (~ n3714) ) ;
 assign n3715 = ( (~ Ng2175)  &  (~ Ng2879) ) | ( (~ Ng2175)  &  (~ Ng2969) ) | ( Ng2879  &  (~ Ng2969) ) ;
 assign Ng20582 = ( (~ n3715) ) ;
 assign n3716 = ( (~ Ng2170)  &  (~ Ng2879) ) | ( (~ Ng2170)  &  (~ Ng2966) ) | ( Ng2879  &  (~ Ng2966) ) ;
 assign Ng20581 = ( (~ n3716) ) ;
 assign n3717 = ( (~ Ng2165)  &  (~ Ng2879) ) | ( (~ Ng2165)  &  (~ Ng2963) ) | ( Ng2879  &  (~ Ng2963) ) ;
 assign Ng20580 = ( (~ n3717) ) ;
 assign n3718 = ( (~ Ng1471)  &  (~ Ng2879) ) | ( (~ Ng1471)  &  (~ Ng2935) ) | ( Ng2879  &  (~ Ng2935) ) ;
 assign Ng20579 = ( (~ n3718) ) ;
 assign n3719 = ( (~ Ng1476)  &  (~ Ng2879) ) | ( (~ Ng1476)  &  (~ Ng2938) ) | ( Ng2879  &  (~ Ng2938) ) ;
 assign Ng20578 = ( (~ n3719) ) ;
 assign n3720 = ( (~ Ng1481)  &  (~ Ng2879) ) | ( (~ Ng1481)  &  (~ Ng2941) ) | ( Ng2879  &  (~ Ng2941) ) ;
 assign Ng20577 = ( (~ n3720) ) ;
 assign n3721 = ( (~ Ng1486)  &  (~ Ng2879) ) | ( (~ Ng1486)  &  (~ Ng2944) ) | ( Ng2879  &  (~ Ng2944) ) ;
 assign Ng20576 = ( (~ n3721) ) ;
 assign n3722 = ( (~ Ng1491)  &  (~ Ng2879) ) | ( (~ Ng1491)  &  (~ Ng2947) ) | ( Ng2879  &  (~ Ng2947) ) ;
 assign Ng20575 = ( (~ n3722) ) ;
 assign n3723 = ( (~ Ng1496)  &  (~ Ng2879) ) | ( (~ Ng1496)  &  (~ Ng2953) ) | ( Ng2879  &  (~ Ng2953) ) ;
 assign Ng20574 = ( (~ n3723) ) ;
 assign n3724 = ( (~ Ng1501)  &  (~ Ng2879) ) | ( (~ Ng1501)  &  (~ Ng2956) ) | ( Ng2879  &  (~ Ng2956) ) ;
 assign Ng20573 = ( (~ n3724) ) ;
 assign n3725 = ( (~ Ng1506)  &  (~ Ng2879) ) | ( (~ Ng1506)  &  (~ Ng2959) ) | ( Ng2879  &  (~ Ng2959) ) ;
 assign Ng20572 = ( (~ n3725) ) ;
 assign n3726 = ( Ng1315  &  (~ Ng2584) ) | ( (~ Ng1315)  &  (~ Ng2704) ) | ( (~ Ng2584)  &  (~ Ng2704) ) ;
 assign Ng20570 = ( (~ n3726) ) ;
 assign n3727 = ( (~ Ng1315)  &  (~ Ng2584) ) | ( Ng1315  &  (~ Ng2631) ) | ( (~ Ng2584)  &  (~ Ng2631) ) ;
 assign Ng20569 = ( (~ n3727) ) ;
 assign n3728 = ( (~ Ng1315)  &  (~ Ng2631) ) | ( Ng1315  &  Ng2628 ) | ( (~ Ng2631)  &  Ng2628 ) ;
 assign Ng20568 = ( (~ n3728) ) ;
 assign n3729 = ( Ng1315  &  (~ Ng1890) ) | ( (~ Ng1315)  &  (~ Ng2010) ) | ( (~ Ng1890)  &  (~ Ng2010) ) ;
 assign Ng20566 = ( (~ n3729) ) ;
 assign n3730 = ( (~ Ng1315)  &  (~ Ng1890) ) | ( Ng1315  &  (~ Ng1937) ) | ( (~ Ng1890)  &  (~ Ng1937) ) ;
 assign Ng20565 = ( (~ n3730) ) ;
 assign n3731 = ( (~ Ng1315)  &  (~ Ng1937) ) | ( Ng1315  &  Ng1934 ) | ( (~ Ng1937)  &  Ng1934 ) ;
 assign Ng20564 = ( (~ n3731) ) ;
 assign n3732 = ( Ng1315  &  (~ Ng1196) ) | ( (~ Ng1315)  &  (~ Ng1316) ) | ( (~ Ng1196)  &  (~ Ng1316) ) ;
 assign Ng20562 = ( (~ n3732) ) ;
 assign n3733 = ( (~ Ng1315)  &  (~ Ng1196) ) | ( Ng1315  &  (~ Ng1243) ) | ( (~ Ng1196)  &  (~ Ng1243) ) ;
 assign Ng20561 = ( (~ n3733) ) ;
 assign n3734 = ( (~ Ng1315)  &  (~ Ng1243) ) | ( Ng1315  &  Ng1240 ) | ( (~ Ng1243)  &  Ng1240 ) ;
 assign Ng20560 = ( (~ n3734) ) ;
 assign n3735 = ( Ng1315  &  (~ Ng510) ) | ( (~ Ng1315)  &  (~ Ng630) ) | ( (~ Ng510)  &  (~ Ng630) ) ;
 assign Ng20558 = ( (~ n3735) ) ;
 assign n3736 = ( (~ Ng1315)  &  (~ Ng510) ) | ( Ng1315  &  (~ Ng557) ) | ( (~ Ng510)  &  (~ Ng557) ) ;
 assign Ng20557 = ( (~ n3736) ) ;
 assign n3737 = ( (~ Ng1315)  &  (~ Ng557) ) | ( Ng1315  &  Ng554 ) | ( (~ Ng557)  &  Ng554 ) ;
 assign Ng20556 = ( (~ n3737) ) ;
 assign n3738 = ( n649 ) | ( n1532 ) ;
 assign n3739 = ( n654 ) | ( n1487 ) ;
 assign n3740 = ( (~ n564)  &  n1300 ) ;
 assign n3741 = ( n659 ) | ( (~ n1300) ) ;
 assign n3742 = ( (~ n569)  &  n1276 ) ;
 assign n3743 = ( n662 ) | ( (~ n1276) ) ;
 assign n3744 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ Ng1315)  &  Ng2812 ) | ( (~ wire1605)  &  Ng2811 ) | ( Ng2812  &  Ng2811 ) ;
 assign n3746 = ( n532  &  (~ n3744) ) | ( wire1603  &  n532  &  (~ Ng2813) ) ;
 assign n3748 = ( Ng2611  &  n679 ) | ( n2278  &  n679 ) | ( Ng2611  &  n1093 ) | ( n2278  &  n1093 ) ;
 assign n3749 = ( n679  &  n2278 ) | ( (~ n1111)  &  n2278 ) | ( n679  &  Ng2610 ) | ( (~ n1111)  &  Ng2610 ) ;
 assign n3750 = ( n679  &  n2278 ) | ( (~ n1106)  &  n2278 ) | ( n679  &  Ng2608 ) | ( (~ n1106)  &  Ng2608 ) ;
 assign n3751 = ( n679  &  n2278 ) | ( (~ n1103)  &  n2278 ) | ( n679  &  Ng2607 ) | ( (~ n1103)  &  Ng2607 ) ;
 assign n3752 = ( n679  &  n2278 ) | ( (~ n1096)  &  n2278 ) | ( n679  &  Ng2606 ) | ( (~ n1096)  &  Ng2606 ) ;
 assign n3754 = ( n679  &  n2278 ) | ( (~ n1109)  &  n2278 ) | ( n679  &  Ng2605 ) | ( (~ n1109)  &  Ng2605 ) ;
 assign n3755 = ( n679  &  n2278 ) | ( (~ n1101)  &  n2278 ) | ( n679  &  Ng2604 ) | ( (~ n1101)  &  Ng2604 ) ;
 assign n3756 = ( n679  &  n2278 ) | ( (~ n1099)  &  n2278 ) | ( n679  &  Ng2603 ) | ( (~ n1099)  &  Ng2603 ) ;
 assign n3758 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ Ng1315)  &  Ng2118 ) | ( (~ wire1605)  &  Ng2117 ) | ( Ng2118  &  Ng2117 ) ;
 assign n3760 = ( n519  &  (~ n3758) ) | ( wire1603  &  n519  &  (~ Ng2119) ) ;
 assign n3762 = ( n675  &  n2291 ) | ( (~ n1087)  &  n2291 ) | ( n675  &  Ng1917 ) | ( (~ n1087)  &  Ng1917 ) ;
 assign n3763 = ( n675  &  n2291 ) | ( (~ n1085)  &  n2291 ) | ( n675  &  Ng1916 ) | ( (~ n1085)  &  Ng1916 ) ;
 assign n3764 = ( n675  &  n2291 ) | ( (~ n1080)  &  n2291 ) | ( n675  &  Ng1914 ) | ( (~ n1080)  &  Ng1914 ) ;
 assign n3765 = ( n675  &  n2291 ) | ( (~ n1077)  &  n2291 ) | ( n675  &  Ng1913 ) | ( (~ n1077)  &  Ng1913 ) ;
 assign n3766 = ( n675  &  n2291 ) | ( (~ n1070)  &  n2291 ) | ( n675  &  Ng1912 ) | ( (~ n1070)  &  Ng1912 ) ;
 assign n3768 = ( n675  &  n2291 ) | ( (~ n1083)  &  n2291 ) | ( n675  &  Ng1911 ) | ( (~ n1083)  &  Ng1911 ) ;
 assign n3769 = ( n675  &  n2291 ) | ( (~ n1075)  &  n2291 ) | ( n675  &  Ng1910 ) | ( (~ n1075)  &  Ng1910 ) ;
 assign n3770 = ( n675  &  n2291 ) | ( (~ n1073)  &  n2291 ) | ( n675  &  Ng1909 ) | ( (~ n1073)  &  Ng1909 ) ;
 assign n3772 = ( n1996  &  n1998 ) | ( n1334  &  n1998 ) | ( n1996  &  n2000 ) | ( n1334  &  n2000 ) ;
 assign n3774 = ( n2000  &  n1996 ) | ( n1334  &  n1996 ) | ( n2000  &  n2002 ) | ( n1334  &  n2002 ) ;
 assign n3776 = ( (~ n1998)  &  (~ n2002) ) | ( (~ n1998)  &  (~ n3772) ) | ( (~ n2002)  &  (~ n3774) ) | ( (~ n3772)  &  (~ n3774) ) ;
 assign n3779 = ( n1325  &  (~ n2005) ) | ( n2003  &  (~ n2005) ) | ( n1325  &  n2006 ) | ( n2003  &  n2006 ) ;
 assign n3781 = ( n1325  &  n2003 ) | ( n2006  &  n2003 ) | ( n1325  &  n2008 ) | ( n2006  &  n2008 ) ;
 assign n3783 = ( n2005  &  (~ n2008) ) | ( n2005  &  (~ n3779) ) | ( (~ n2008)  &  (~ n3781) ) | ( (~ n3779)  &  (~ n3781) ) ;
 assign n3785 = ( n2029  &  n2031 ) | ( n1367  &  n2031 ) | ( n2029  &  n2033 ) | ( n1367  &  n2033 ) ;
 assign n3787 = ( n2033  &  n2029 ) | ( n1367  &  n2029 ) | ( n2033  &  n2035 ) | ( n1367  &  n2035 ) ;
 assign n3789 = ( (~ n2031)  &  (~ n2035) ) | ( (~ n2031)  &  (~ n3785) ) | ( (~ n2035)  &  (~ n3787) ) | ( (~ n3785)  &  (~ n3787) ) ;
 assign n3792 = ( n1358  &  (~ n2038) ) | ( n2036  &  (~ n2038) ) | ( n1358  &  n2039 ) | ( n2036  &  n2039 ) ;
 assign n3794 = ( n1358  &  n2036 ) | ( n2039  &  n2036 ) | ( n1358  &  n2041 ) | ( n2039  &  n2041 ) ;
 assign n3796 = ( n2038  &  (~ n2041) ) | ( n2038  &  (~ n3792) ) | ( (~ n2041)  &  (~ n3794) ) | ( (~ n3792)  &  (~ n3794) ) ;
 assign n3798 = ( n2062  &  n2064 ) | ( n1400  &  n2064 ) | ( n2062  &  n2066 ) | ( n1400  &  n2066 ) ;
 assign n3800 = ( n2066  &  n2062 ) | ( n1400  &  n2062 ) | ( n2066  &  n2068 ) | ( n1400  &  n2068 ) ;
 assign n3802 = ( (~ n2064)  &  (~ n2068) ) | ( (~ n2064)  &  (~ n3798) ) | ( (~ n2068)  &  (~ n3800) ) | ( (~ n3798)  &  (~ n3800) ) ;
 assign n3805 = ( n1391  &  (~ n2071) ) | ( n2069  &  (~ n2071) ) | ( n1391  &  n2072 ) | ( n2069  &  n2072 ) ;
 assign n3807 = ( n1391  &  n2069 ) | ( n2072  &  n2069 ) | ( n1391  &  n2074 ) | ( n2072  &  n2074 ) ;
 assign n3809 = ( n2071  &  (~ n2074) ) | ( n2071  &  (~ n3805) ) | ( (~ n2074)  &  (~ n3807) ) | ( (~ n3805)  &  (~ n3807) ) ;
 assign n3811 = ( n2095  &  n2097 ) | ( n1433  &  n2097 ) | ( n2095  &  n2099 ) | ( n1433  &  n2099 ) ;
 assign n3813 = ( n2099  &  n2095 ) | ( n1433  &  n2095 ) | ( n2099  &  n2101 ) | ( n1433  &  n2101 ) ;
 assign n3815 = ( (~ n2097)  &  (~ n2101) ) | ( (~ n2097)  &  (~ n3811) ) | ( (~ n2101)  &  (~ n3813) ) | ( (~ n3811)  &  (~ n3813) ) ;
 assign n3818 = ( n1424  &  (~ n2104) ) | ( n2102  &  (~ n2104) ) | ( n1424  &  n2105 ) | ( n2102  &  n2105 ) ;
 assign n3820 = ( n1424  &  n2102 ) | ( n2105  &  n2102 ) | ( n1424  &  n2107 ) | ( n2105  &  n2107 ) ;
 assign n3822 = ( n2104  &  (~ n2107) ) | ( n2104  &  (~ n3818) ) | ( (~ n2107)  &  (~ n3820) ) | ( (~ n3818)  &  (~ n3820) ) ;
 assign n3824 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ Ng1315)  &  Ng1424 ) | ( (~ wire1605)  &  Ng1423 ) | ( Ng1424  &  Ng1423 ) ;
 assign n3826 = ( n433 ) | ( n358 ) | ( n515 ) | ( n282 ) | ( n256 ) | ( n317 ) ;
 assign n3828 = ( n671  &  n2444 ) | ( (~ n1034)  &  n2444 ) | ( n671  &  Ng1223 ) | ( (~ n1034)  &  Ng1223 ) ;
 assign n3829 = ( n671  &  n2444 ) | ( (~ n1032)  &  n2444 ) | ( n671  &  Ng1222 ) | ( (~ n1032)  &  Ng1222 ) ;
 assign n3830 = ( n671  &  n2444 ) | ( (~ n1027)  &  n2444 ) | ( n671  &  Ng1220 ) | ( (~ n1027)  &  Ng1220 ) ;
 assign n3831 = ( n671  &  n2444 ) | ( (~ n1024)  &  n2444 ) | ( n671  &  Ng1219 ) | ( (~ n1024)  &  Ng1219 ) ;
 assign n3832 = ( n671  &  n2444 ) | ( (~ n1036)  &  n2444 ) | ( n671  &  Ng1218 ) | ( (~ n1036)  &  Ng1218 ) ;
 assign n3833 = ( n671  &  n2444 ) | ( (~ n1030)  &  n2444 ) | ( n671  &  Ng1217 ) | ( (~ n1030)  &  Ng1217 ) ;
 assign n3834 = ( n671  &  n2444 ) | ( (~ n1021)  &  n2444 ) | ( n671  &  Ng1216 ) | ( (~ n1021)  &  Ng1216 ) ;
 assign n3835 = ( n671  &  n2444 ) | ( (~ n1017)  &  n2444 ) | ( n671  &  Ng1215 ) | ( (~ n1017)  &  Ng1215 ) ;
 assign n3836 = ( (~ wire1605)  &  (~ Ng1315) ) | ( (~ Ng1315)  &  Ng738 ) | ( (~ wire1605)  &  Ng737 ) | ( Ng738  &  Ng737 ) ;
 assign n3838 = ( n383 ) | ( n308 ) | ( n493 ) | ( n247 ) | ( n228 ) | ( n275 ) ;
 assign n3840 = ( n667  &  n2467 ) | ( (~ n1007)  &  n2467 ) | ( n667  &  Ng537 ) | ( (~ n1007)  &  Ng537 ) ;
 assign n3841 = ( n667  &  n2467 ) | ( (~ n1005)  &  n2467 ) | ( n667  &  Ng536 ) | ( (~ n1005)  &  Ng536 ) ;
 assign n3842 = ( n667  &  n2467 ) | ( (~ n999)  &  n2467 ) | ( n667  &  Ng534 ) | ( (~ n999)  &  Ng534 ) ;
 assign n3843 = ( n667  &  n2467 ) | ( (~ n996)  &  n2467 ) | ( n667  &  Ng533 ) | ( (~ n996)  &  Ng533 ) ;
 assign n3844 = ( n667  &  n2467 ) | ( (~ n1009)  &  n2467 ) | ( n667  &  Ng532 ) | ( (~ n1009)  &  Ng532 ) ;
 assign n3845 = ( n667  &  n2467 ) | ( (~ n1002)  &  n2467 ) | ( n667  &  Ng531 ) | ( (~ n1002)  &  Ng531 ) ;
 assign n3846 = ( n667  &  n2467 ) | ( (~ n992)  &  n2467 ) | ( n667  &  Ng530 ) | ( (~ n992)  &  Ng530 ) ;
 assign n3847 = ( n667  &  n2467 ) | ( (~ n1011)  &  n2467 ) | ( n667  &  Ng529 ) | ( (~ n1011)  &  Ng529 ) ;
 assign n3849 = ( n94 ) | ( n109 ) | ( n623 ) ;
 assign n3848 = ( n3849  &  n2534 ) | ( n3849  &  n1654 ) ;
 assign n3850 = ( (~ n103)  &  (~ n611) ) | ( (~ n103)  &  n1646 ) | ( (~ n611)  &  n2534 ) | ( n1646  &  n2534 ) ;
 assign n3852 = ( n82 ) | ( n100 ) | ( n609 ) ;
 assign n3851 = ( n3852  &  n2560 ) | ( n3852  &  n1689 ) ;
 assign n3853 = ( (~ n91)  &  (~ n597) ) | ( (~ n91)  &  n1681 ) | ( (~ n597)  &  n2560 ) | ( n1681  &  n2560 ) ;
 assign n3855 = ( n73 ) | ( n88 ) | ( n595 ) ;
 assign n3854 = ( n3855  &  n2584 ) | ( n3855  &  n1724 ) ;
 assign n3856 = ( (~ n79)  &  (~ n583) ) | ( (~ n79)  &  n1716 ) | ( (~ n583)  &  n2584 ) | ( n1716  &  n2584 ) ;
 assign n3858 = ( n66 ) | ( n76 ) | ( n581 ) ;
 assign n3857 = ( n3858  &  n2608 ) | ( n3858  &  n1759 ) ;
 assign n3859 = ( (~ n70)  &  (~ n574) ) | ( (~ n70)  &  n1751 ) | ( (~ n574)  &  n2608 ) | ( n1751  &  n2608 ) ;
 assign n3860 = ( n2497 ) | ( (~ n4456) ) ;
 assign n3861 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng2253 ) | ( (~ Ng853)  &  Ng2254 ) | ( Ng2253  &  Ng2254 ) ;
 assign n3862 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng1559 ) | ( (~ Ng853)  &  Ng1560 ) | ( Ng1559  &  Ng1560 ) ;
 assign n3863 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng865 ) | ( (~ Ng853)  &  Ng866 ) | ( Ng865  &  Ng866 ) ;
 assign n3864 = ( (~ wire1612)  &  (~ Ng853) ) | ( (~ wire1612)  &  Ng177 ) | ( (~ Ng853)  &  Ng178 ) | ( Ng177  &  Ng178 ) ;
 assign n3869 = ( n2189 ) | ( n2191 ) | ( n2192 ) ;
 assign n3870 = ( n2198 ) | ( n2199 ) | ( n2201 ) | ( n2203 ) | ( n2204 ) | ( n2194 ) | ( n2196 ) | ( n3869 ) ;
 assign n3871 = ( (~ Ng1315) ) | ( Ng2802 ) ;
 assign n3872 = ( n2205 ) | ( n2207 ) | ( n2208 ) ;
 assign n3873 = ( n2214 ) | ( n2215 ) | ( n2217 ) | ( n2219 ) | ( n2220 ) | ( n2210 ) | ( n2212 ) | ( n3872 ) ;
 assign n3874 = ( (~ Ng1315) ) | ( Ng2108 ) ;
 assign n3875 = ( n2221 ) | ( n2223 ) | ( n2225 ) ;
 assign n3876 = ( n2231 ) | ( n2233 ) | ( n2235 ) | ( n2237 ) | ( n2239 ) | ( n2227 ) | ( n2229 ) | ( n3875 ) ;
 assign n3877 = ( (~ Ng1315) ) | ( Ng1414 ) ;
 assign n3878 = ( n2241 ) | ( n2243 ) | ( n2245 ) ;
 assign n3879 = ( n2251 ) | ( n2253 ) | ( n2255 ) | ( n2257 ) | ( n2259 ) | ( n2247 ) | ( n2249 ) | ( n3878 ) ;
 assign n3880 = ( (~ Ng1315) ) | ( Ng728 ) ;
 assign n3881 = ( Ng3139  &  n2453 ) | ( n2453  &  (~ n4878) ) ;
 assign n3884 = ( wire1605 ) | ( Ng8284 ) | ( (~ Ng548) ) ;
 assign n3886 = ( wire1605  &  n2727 ) | ( (~ wire1605)  &  (~ Ng1234) ) | ( n2727  &  (~ Ng1234) ) ;
 assign n3889 = ( wire1605  &  n2728 ) | ( (~ wire1605)  &  (~ Ng1928) ) | ( n2728  &  (~ Ng1928) ) ;
 assign n3892 = ( wire1605  &  n2729 ) | ( (~ wire1605)  &  (~ Ng2622) ) | ( n2729  &  (~ Ng2622) ) ;
 assign n3895 = ( n331  &  n569 ) | ( (~ n331)  &  n3742 ) | ( n569  &  n3742 ) ;
 assign n3897 = ( Pg3229  &  Ng2612 ) | ( (~ Pg3229)  &  Ng2615 ) | ( Ng2612  &  Ng2615 ) ;
 assign n3898 = ( n1191  &  n1193 ) | ( (~ n1191)  &  (~ n1193) ) ;
 assign n3900 = ( Ng2631 ) | ( n2278 ) | ( (~ n3897) ) ;
 assign n3904 = ( Pg3229  &  Ng1918 ) | ( (~ Pg3229)  &  Ng1921 ) | ( Ng1918  &  Ng1921 ) ;
 assign n3905 = ( n1177  &  n1179 ) | ( (~ n1177)  &  (~ n1179) ) ;
 assign n3907 = ( Ng1937 ) | ( n2291 ) | ( (~ n3904) ) ;
 assign n3909 = ( (~ n567)  &  n2324 ) | ( (~ n177)  &  (~ n567)  &  (~ n1545) ) ;
 assign n3910 = ( n562  &  n3909 ) | ( n562  &  n567  &  (~ n1966) ) ;
 assign n3912 = ( n555  &  (~ n562) ) | ( (~ n562)  &  n1067 ) ;
 assign n3913 = ( (~ n555)  &  n562  &  (~ n1067) ) | ( n562  &  n567  &  (~ n1067) ) ;
 assign n3916 = ( (~ n923) ) | ( n3912 ) | ( n3913 ) ;
 assign n3925 = ( (~ n560)  &  n2359 ) | ( (~ n173)  &  (~ n560)  &  (~ n1555) ) ;
 assign n3926 = ( n553  &  n3925 ) | ( n553  &  n560  &  (~ n1968) ) ;
 assign n3928 = ( n546  &  (~ n553) ) | ( (~ n553)  &  n1064 ) ;
 assign n3929 = ( (~ n546)  &  n553  &  (~ n1064) ) | ( n553  &  n560  &  (~ n1064) ) ;
 assign n3932 = ( (~ n918) ) | ( n3928 ) | ( n3929 ) ;
 assign n3941 = ( (~ n551)  &  n2394 ) | ( (~ n167)  &  (~ n551)  &  (~ n1565) ) ;
 assign n3942 = ( n544  &  n3941 ) | ( n544  &  n551  &  (~ n1970) ) ;
 assign n3944 = ( n540  &  (~ n544) ) | ( (~ n544)  &  n1061 ) ;
 assign n3945 = ( (~ n540)  &  n544  &  (~ n1061) ) | ( n544  &  n551  &  (~ n1061) ) ;
 assign n3948 = ( (~ n913) ) | ( n3944 ) | ( n3945 ) ;
 assign n3957 = ( (~ n542)  &  n2429 ) | ( (~ n160)  &  (~ n542)  &  (~ n1575) ) ;
 assign n3958 = ( n538  &  n3957 ) | ( n538  &  n542  &  (~ n1972) ) ;
 assign n3960 = ( n534  &  (~ n538) ) | ( (~ n538)  &  n1058 ) ;
 assign n3961 = ( (~ n534)  &  n538  &  (~ n1058) ) | ( n538  &  n542  &  (~ n1058) ) ;
 assign n3964 = ( (~ n908) ) | ( n3960 ) | ( n3961 ) ;
 assign n3973 = ( n562  &  (~ n567) ) | ( n562  &  (~ Ng2257) ) | ( n562  &  n2320 ) ;
 assign n3978 = ( n553  &  (~ n560) ) | ( n553  &  (~ Ng2257) ) | ( n553  &  n2355 ) ;
 assign n3983 = ( n544  &  (~ n551) ) | ( n544  &  (~ Ng2257) ) | ( n544  &  n2390 ) ;
 assign n3988 = ( n538  &  (~ n542) ) | ( n538  &  (~ Ng2257) ) | ( n538  &  n2425 ) ;
 assign n3993 = ( n450  &  n1458 ) | ( (~ n450)  &  (~ n1458) ) ;
 assign n3994 = ( n265  &  n1455 ) | ( (~ n265)  &  (~ n1455) ) ;
 assign n3996 = ( n2327 ) | ( n2020 ) | ( n521 ) ;
 assign n3995 = ( (~ n521)  &  n3996 ) | ( (~ n2020)  &  (~ n2327)  &  n3996 ) ;
 assign n3997 = ( n400  &  n1466 ) | ( (~ n400)  &  (~ n1466) ) ;
 assign n3998 = ( n237  &  n1463 ) | ( (~ n237)  &  (~ n1463) ) ;
 assign n4000 = ( n2362 ) | ( n2053 ) | ( n499 ) ;
 assign n3999 = ( (~ n499)  &  n4000 ) | ( (~ n2053)  &  (~ n2362)  &  n4000 ) ;
 assign n4001 = ( n350  &  n1474 ) | ( (~ n350)  &  (~ n1474) ) ;
 assign n4002 = ( n214  &  n1471 ) | ( (~ n214)  &  (~ n1471) ) ;
 assign n4004 = ( n2397 ) | ( n2086 ) | ( n464 ) ;
 assign n4003 = ( (~ n464)  &  n4004 ) | ( (~ n2086)  &  (~ n2397)  &  n4004 ) ;
 assign n4005 = ( n300  &  n1482 ) | ( (~ n300)  &  (~ n1482) ) ;
 assign n4006 = ( n197  &  n1479 ) | ( (~ n197)  &  (~ n1479) ) ;
 assign n4008 = ( n2432 ) | ( n2119 ) | ( n419 ) ;
 assign n4007 = ( (~ n419)  &  n4008 ) | ( (~ n2119)  &  (~ n2432)  &  n4008 ) ;
 assign n4010 = ( wire1603 ) | ( Pg16297 ) | ( Ng506 ) ;
 assign Ng23154 = ( (~ Ng506)  &  n4010 ) | ( n4010  &  Ng507 ) ;
 assign n4011 = ( Pg16355  &  (~ wire1603) ) | ( Pg16355  &  Ng23154 ) | ( wire1603  &  Ng23154 ) ;
 assign Ng27212 = ( n4011  &  (~ Ng1192) ) | ( n4011  &  Ng1193 ) | ( Ng1192  &  Ng1193 ) ;
 assign n4013 = ( Pg16399  &  (~ wire1603) ) | ( Pg16399  &  Ng27212 ) | ( wire1603  &  Ng27212 ) ;
 assign n4016 = ( (~ Pg16437)  &  (~ wire1603) ) | ( (~ Pg16437)  &  (~ Ng29440) ) | ( wire1603  &  (~ Ng29440) ) ;
 assign n4020 = ( Ng298 ) | ( Ng299 ) ;
 assign n4022 = ( wire1594  &  n2929 ) | ( (~ wire1594)  &  (~ Ng992) ) | ( n2929  &  (~ Ng992) ) ;
 assign n4025 = ( wire1594  &  n2930 ) | ( (~ wire1594)  &  (~ Ng1686) ) | ( n2930  &  (~ Ng1686) ) ;
 assign n4028 = ( wire1594  &  n2931 ) | ( (~ wire1594)  &  (~ Ng2380) ) | ( n2931  &  (~ Ng2380) ) ;
 assign n4031 = ( Pg3229  &  Ng1224 ) | ( (~ Pg3229)  &  Ng1227 ) | ( Ng1224  &  Ng1227 ) ;
 assign n4032 = ( n1163  &  n1165 ) | ( (~ n1163)  &  (~ n1165) ) ;
 assign n4034 = ( Ng1243 ) | ( n2444 ) | ( (~ n4031) ) ;
 assign n4037 = ( (~ n923) ) | ( n1507 ) ;
 assign n4041 = ( (~ n918) ) | ( n1511 ) ;
 assign n4045 = ( (~ n913) ) | ( n1515 ) ;
 assign n4049 = ( (~ n908) ) | ( n1519 ) ;
 assign n4054 = ( Pg3229  &  Ng538 ) | ( (~ Pg3229)  &  Ng541 ) | ( Ng538  &  Ng541 ) ;
 assign n4055 = ( n1149  &  n1151 ) | ( (~ n1149)  &  (~ n1151) ) ;
 assign n4057 = ( Ng557 ) | ( n2467 ) | ( (~ n4054) ) ;
 assign n4059 = ( n629  &  n1537 ) | ( (~ n629)  &  (~ n1537) ) ;
 assign n4060 = ( (~ n1546)  &  Ng2257 ) | ( n1546  &  n2323 ) | ( Ng2257  &  n2323 ) ;
 assign n4062 = ( Ng853  &  n4060 ) ;
 assign n4066 = ( wire1594  &  n4060 ) ;
 assign n4069 = ( wire1612  &  n4060 ) ;
 assign n4071 = ( n615  &  n1547 ) | ( (~ n615)  &  (~ n1547) ) ;
 assign n4072 = ( (~ n1556)  &  Ng2257 ) | ( n1556  &  n2358 ) | ( Ng2257  &  n2358 ) ;
 assign n4074 = ( Ng853  &  n4072 ) ;
 assign n4078 = ( wire1594  &  n4072 ) ;
 assign n4081 = ( wire1612  &  n4072 ) ;
 assign n4083 = ( n601  &  n1557 ) | ( (~ n601)  &  (~ n1557) ) ;
 assign n4084 = ( (~ n1566)  &  Ng2257 ) | ( n1566  &  n2393 ) | ( Ng2257  &  n2393 ) ;
 assign n4086 = ( Ng853  &  n4084 ) ;
 assign n4090 = ( wire1594  &  n4084 ) ;
 assign n4093 = ( wire1612  &  n4084 ) ;
 assign n4095 = ( n587  &  n1567 ) | ( (~ n587)  &  (~ n1567) ) ;
 assign n4096 = ( (~ n1576)  &  Ng2257 ) | ( n1576  &  n2428 ) | ( Ng2257  &  n2428 ) ;
 assign n4098 = ( Ng853  &  n4096 ) ;
 assign n4102 = ( wire1594  &  n4096 ) ;
 assign n4105 = ( wire1612  &  n4096 ) ;
 assign n4108 = ( n1593 ) | ( n891 ) ;
 assign n4107 = ( (~ n620)  &  n4108 ) | ( n620  &  (~ n4108) ) ;
 assign n4110 = ( n1600 ) | ( n887 ) ;
 assign n4109 = ( (~ n606)  &  n4110 ) | ( n606  &  (~ n4110) ) ;
 assign n4112 = ( n1607 ) | ( n883 ) ;
 assign n4111 = ( (~ n592)  &  n4112 ) | ( n592  &  (~ n4112) ) ;
 assign n4114 = ( n1614 ) | ( n880 ) ;
 assign n4113 = ( (~ n578)  &  n4114 ) | ( n578  &  (~ n4114) ) ;
 assign n4118 = ( n2547 ) | ( n569 ) ;
 assign n4116 = ( n2545  &  n4118 ) | ( (~ n2547)  &  n4118 ) | ( (~ n3003)  &  n4118 ) ;
 assign n4120 = ( n662  &  (~ n2547) ) | ( n662  &  (~ n3007) ) | ( n2547  &  (~ n3007) ) ;
 assign n4123 = ( n2547 ) | ( n564 ) ;
 assign n4122 = ( (~ n2547)  &  n4123 ) | ( n2571  &  n4123 ) | ( (~ n3016)  &  n4123 ) ;
 assign n4125 = ( n659  &  (~ n2547) ) | ( n659  &  (~ n3020) ) | ( n2547  &  (~ n3020) ) ;
 assign n4128 = ( n2547 ) | ( n557 ) ;
 assign n4127 = ( (~ n2547)  &  n4128 ) | ( n2595  &  n4128 ) | ( (~ n3029)  &  n4128 ) ;
 assign n4130 = ( n654  &  (~ n2547) ) | ( n654  &  (~ n3033) ) | ( n2547  &  (~ n3033) ) ;
 assign n4133 = ( n2547 ) | ( n548 ) ;
 assign n4132 = ( (~ n2547)  &  n4133 ) | ( n2619  &  n4133 ) | ( (~ n3042)  &  n4133 ) ;
 assign n4135 = ( n649  &  (~ n2547) ) | ( n649  &  (~ n3046) ) | ( n2547  &  (~ n3046) ) ;
 assign n4136 = ( (~ n455) ) | ( n488 ) | ( n1786 ) ;
 assign n4137 = ( (~ n405) ) | ( n443 ) | ( n1797 ) ;
 assign n4138 = ( (~ n355) ) | ( n393 ) | ( n1807 ) ;
 assign n4139 = ( (~ n305) ) | ( n343 ) | ( n1817 ) ;
 assign n4140 = ( (~ Ng1315) ) | ( n745 ) ;
 assign n4142 = ( n1640  &  n4150 ) ;
 assign n4144 = ( (~ wire1603) ) | ( n745 ) ;
 assign n4147 = ( (~ wire1605) ) | ( n745 ) ;
 assign n4150 = ( Pg3229  &  n599 ) | ( (~ Pg3229)  &  (~ n599) ) ;
 assign n4158 = ( (~ n599)  &  n611  &  n632 ) | ( (~ n599)  &  (~ n623)  &  n632 ) ;
 assign n4163 = ( Ng853  &  n731 ) ;
 assign n4165 = ( n509  &  n2138  &  n486 ) ;
 assign n4167 = ( wire1594  &  n731 ) ;
 assign n4170 = ( wire1612  &  n731 ) ;
 assign n4181 = ( (~ n453)  &  n486  &  n524 ) | ( (~ n453)  &  (~ n509)  &  n524 ) ;
 assign n4187 = ( (~ Ng1315) ) | ( n740 ) ;
 assign n4189 = ( n1675  &  n4197 ) ;
 assign n4191 = ( (~ wire1603) ) | ( n740 ) ;
 assign n4194 = ( (~ wire1605) ) | ( n740 ) ;
 assign n4197 = ( Pg3229  &  n585 ) | ( (~ Pg3229)  &  (~ n585) ) ;
 assign n4205 = ( (~ n585)  &  n597  &  n618 ) | ( (~ n585)  &  (~ n609)  &  n618 ) ;
 assign n4210 = ( Ng853  &  n728 ) ;
 assign n4212 = ( n474  &  n2139  &  n441 ) ;
 assign n4214 = ( wire1594  &  n728 ) ;
 assign n4217 = ( wire1612  &  n728 ) ;
 assign n4228 = ( (~ n403)  &  n441  &  n502 ) | ( (~ n403)  &  (~ n474)  &  n502 ) ;
 assign n4234 = ( (~ Ng1315) ) | ( n739 ) ;
 assign n4236 = ( n1710  &  n4244 ) ;
 assign n4238 = ( (~ wire1603) ) | ( n739 ) ;
 assign n4241 = ( (~ wire1605) ) | ( n739 ) ;
 assign n4244 = ( Pg3229  &  n576 ) | ( (~ Pg3229)  &  (~ n576) ) ;
 assign n4252 = ( (~ n576)  &  n583  &  n604 ) | ( (~ n576)  &  (~ n595)  &  n604 ) ;
 assign n4257 = ( Ng853  &  n724 ) ;
 assign n4259 = ( n429  &  n2140  &  n391 ) ;
 assign n4261 = ( wire1594  &  n724 ) ;
 assign n4264 = ( wire1612  &  n724 ) ;
 assign n4275 = ( (~ n353)  &  n391  &  n467 ) | ( (~ n353)  &  (~ n429)  &  n467 ) ;
 assign n4281 = ( (~ Ng1315) ) | ( n736 ) ;
 assign n4283 = ( n1745  &  n4291 ) ;
 assign n4285 = ( (~ wire1603) ) | ( n736 ) ;
 assign n4288 = ( (~ wire1605) ) | ( n736 ) ;
 assign n4291 = ( Pg3229  &  n572 ) | ( (~ Pg3229)  &  (~ n572) ) ;
 assign n4299 = ( (~ n572)  &  n574  &  n590 ) | ( (~ n572)  &  (~ n581)  &  n590 ) ;
 assign n4304 = ( Ng853  &  n719 ) ;
 assign n4306 = ( n379  &  n2141  &  n341 ) ;
 assign n4308 = ( wire1594  &  n719 ) ;
 assign n4311 = ( wire1612  &  n719 ) ;
 assign n4322 = ( (~ n303)  &  n341  &  n422 ) | ( (~ n303)  &  (~ n379)  &  n422 ) ;
 assign n4328 = ( n488  &  n4873 ) | ( (~ n488)  &  (~ n4873) ) ;
 assign n4329 = ( n455  &  n4893 ) | ( (~ n455)  &  (~ n4893) ) ;
 assign n4330 = ( n443  &  n4872 ) | ( (~ n443)  &  (~ n4872) ) ;
 assign n4331 = ( n405  &  n4894 ) | ( (~ n405)  &  (~ n4894) ) ;
 assign n4332 = ( n393  &  n4871 ) | ( (~ n393)  &  (~ n4871) ) ;
 assign n4333 = ( n355  &  n4895 ) | ( (~ n355)  &  (~ n4895) ) ;
 assign n4334 = ( n343  &  n4870 ) | ( (~ n343)  &  (~ n4870) ) ;
 assign n4335 = ( n305  &  n4896 ) | ( (~ n305)  &  (~ n4896) ) ;
 assign n4336 = ( (~ n124) ) | ( (~ n569) ) | ( (~ Ng2584) ) ;
 assign n4337 = ( (~ Ng853) ) | ( (~ Ng2257) ) ;
 assign n4339 = ( n153  &  (~ n1545) ) ;
 assign n4341 = ( (~ wire1594) ) | ( (~ Ng2257) ) ;
 assign n4344 = ( (~ wire1612) ) | ( (~ Ng2257) ) ;
 assign n4347 = ( (~ n121) ) | ( (~ n564) ) | ( (~ Ng1890) ) ;
 assign n4349 = ( n144  &  (~ n1555) ) ;
 assign n4352 = ( (~ n118) ) | ( (~ n557) ) | ( (~ Ng1196) ) ;
 assign n4354 = ( n137  &  (~ n1565) ) ;
 assign n4357 = ( (~ n115) ) | ( (~ n548) ) | ( (~ Ng510) ) ;
 assign n4359 = ( n130  &  (~ n1575) ) ;
 assign n4362 = ( Ng13475  &  Ng2993 ) | ( (~ Ng13475)  &  (~ Ng2993) ) ;
 assign n4370 = ( (~ Ng853) ) | ( n2703 ) ;
 assign n4373 = ( (~ wire1594) ) | ( n2703 ) ;
 assign n4375 = ( (~ wire1612) ) | ( n2703 ) ;
 assign n4385 = ( (~ Ng2185) ) | ( Ng2190 ) | ( Ng2195 ) | ( (~ Ng2200) ) ;
 assign n4404 = ( (~ Ng1491) ) | ( Ng1496 ) | ( Ng1501 ) | ( (~ Ng1506) ) ;
 assign n4423 = ( (~ Ng801) ) | ( Ng805 ) | ( Ng809 ) | ( (~ Ng813) ) ;
 assign n4442 = ( (~ Ng113) ) | ( Ng117 ) | ( Ng121 ) | ( (~ Ng125) ) ;
 assign n4445 = ( n2547 ) | ( n1659 ) ;
 assign n4446 = ( n2547 ) | ( n693 ) ;
 assign n4447 = ( n1916  &  n792 ) ;
 assign n4449 = ( n2547 ) | ( n1694 ) ;
 assign n4450 = ( n2547 ) | ( n689 ) ;
 assign n4451 = ( n2547 ) | ( n1729 ) ;
 assign n4452 = ( n2547 ) | ( n685 ) ;
 assign n4453 = ( n2547 ) | ( n1764 ) ;
 assign n4454 = ( n2547 ) | ( n681 ) ;
 assign n4456 = ( Ng2985 ) | ( Ng2984 ) ;
 assign n4455 = ( (~ Ng3147)  &  (~ n3881) ) | ( (~ Ng3147)  &  (~ Ng3120)  &  n4456 ) ;
 assign n4503 = ( (~ wire1594) ) | ( (~ Ng2257) ) ;
 assign n4506 = ( (~ wire1612) ) | ( (~ Ng2257) ) ;
 assign n4644 = ( n2724  &  n4897 ) | ( (~ n2724)  &  (~ n4897) ) ;
 assign n4869 = ( Ng3002 ) | ( Ng3013 ) | ( Ng3024 ) | ( Ng3006 ) | ( Ng3010 ) ;
 assign Ng20567 = ( (~ n2703) ) ;
 assign n4870 = ( n127 ) | ( (~ Ng2257) ) | ( n2680 ) ;
 assign n4871 = ( n135 ) | ( (~ Ng2257) ) | ( n2671 ) ;
 assign n4872 = ( n142 ) | ( (~ Ng2257) ) | ( n2662 ) ;
 assign n4873 = ( n151 ) | ( (~ Ng2257) ) | ( n2653 ) ;
 assign n4878 = ( Ng2991 ) | ( Ng2992 ) ;
 assign n4893 = ( (~ Ng2257) ) | ( n2715 ) ;
 assign n4894 = ( (~ Ng2257) ) | ( n2716 ) ;
 assign n4895 = ( (~ Ng2257) ) | ( n2717 ) ;
 assign n4896 = ( (~ Ng2257) ) | ( n2718 ) ;
 assign n4897 = ( Pg3231 ) | ( (~ Ng3139) ) ;
 assign n4898 = ( Pg3231 ) | ( (~ Ng3120) ) ;
 assign n4900 = ( (~ n2725)  &  n4897 ) | ( n2725  &  (~ n4897) ) ;
 assign n4904 = ( n486  &  n524  &  (~ n2138) ) ;
 assign n4905 = ( n441  &  n502  &  (~ n2139) ) ;
 assign n4906 = ( n391  &  n467  &  (~ n2140) ) ;
 assign n4907 = ( n341  &  n422  &  (~ n2141) ) ;
 assign Pg25442 = ( wire1521 ) ;
 assign Pg25420 = ( wire1521 ) ;
 assign Pg8167 = ( wire1594 ) ;
 assign Pg8106 = ( wire1605 ) ;
 assign Pg8087 = ( wire1612 ) ;
 assign Pg8082 = ( wire1594 ) ;
 assign Pg8030 = ( wire1603 ) ;
 assign Pg8012 = ( wire1612 ) ;
 assign Pg8007 = ( wire1594 ) ;
 assign Pg7961 = ( wire1612 ) ;
 assign Pg7956 = ( wire1594 ) ;
 assign Pg7909 = ( wire1612 ) ;
 assign Pg7487 = ( wire1603 ) ;
 assign Pg7425 = ( wire1605 ) ;
 assign Pg7390 = ( wire1603 ) ;
 assign Pg7357 = ( wire1603 ) ;
 assign Pg7302 = ( wire1605 ) ;
 assign Pg7264 = ( wire1594 ) ;
 assign Pg7229 = ( wire1605 ) ;
 assign Pg7194 = ( wire1603 ) ;
 assign Pg7161 = ( wire1603 ) ;
 assign Pg7084 = ( wire1594 ) ;
 assign Pg7052 = ( wire1605 ) ;
 assign Pg7014 = ( wire1594 ) ;
 assign Pg6979 = ( wire1605 ) ;
 assign Pg6944 = ( wire1603 ) ;
 assign Pg6911 = ( wire1603 ) ;
 assign Pg6837 = ( wire1612 ) ;
 assign Pg6782 = ( wire1594 ) ;
 assign Pg6750 = ( wire1605 ) ;
 assign Pg6712 = ( wire1594 ) ;
 assign Pg6677 = ( wire1605 ) ;
 assign Pg6642 = ( wire1603 ) ;
 assign Pg6573 = ( wire1612 ) ;
 assign Pg6518 = ( wire1594 ) ;
 assign Pg6485 = ( wire1605 ) ;
 assign Pg6447 = ( wire1594 ) ;
 assign Pg6368 = ( wire1612 ) ;
 assign Pg6313 = ( wire1594 ) ;
 assign Pg6231 = ( wire1612 ) ;
 assign Pg5796 = ( wire1603 ) ;
 assign Pg5747 = ( wire1605 ) ;
 assign Pg5738 = ( wire1603 ) ;
 assign Pg5695 = ( wire1605 ) ;
 assign Pg5686 = ( wire1603 ) ;
 assign Pg5657 = ( wire1605 ) ;
 assign Pg5648 = ( wire1603 ) ;
 assign Pg5637 = ( wire1609 ) ;
 assign Pg5629 = ( wire1605 ) ;
 assign Pg5612 = ( wire1609 ) ;
 assign Pg5595 = ( wire1609 ) ;
 assign Pg5555 = ( wire1612 ) ;
 assign Pg5549 = ( wire1609 ) ;
 assign Pg5511 = ( wire1612 ) ;
 assign Pg5472 = ( wire1612 ) ;
 assign Pg5437 = ( wire1612 ) ;


endmodule

