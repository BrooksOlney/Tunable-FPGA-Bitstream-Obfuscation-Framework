// sk = 101111100100001001010
`timescale 10ns/1ns
module apex4 (/* input clk, */ input [20:0] sk, input i_0_, input i_1_, input i_2_, input i_6_, input i_7_, input i_8_, input i_3_, input i_4_, input i_5_, output wire o_1_, output wire o_2_, output wire o_3_, output wire o_4_, output wire o_5_, output wire o_6_, output wire o_7_, output wire o_8_, output wire o_9_, output wire o_10_, output wire o_11_, output wire o_12_, output wire o_13_, output wire o_14_, output wire o_15_, output wire o_16_, output wire o_17_, output wire o_18_);

//reg [8:0] inputs;
//reg [17:0] outputs;
//reg [20:0] sk_reg;
//always @(posedge clk) inputs = {i_0_, i_1_, i_2_, i_6_, i_7_, i_8_, i_3_, i_4_, i_5_};
//always @(posedge clk) outputs = {o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_};
//always @(posedge clk) sk_reg = {o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_, o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_};

	wire g82, g199, g263, g320, g356, g395, g418, g437, g454, g467, g490;
	wire g510, g520, g523, g532, g537, g540, g542, g1, g2, g3, g4;
	wire g5, g6, g7, g8, g9, g10, g11, g12, g13, g14, g15;
	wire g16, g17, g18, g19, g20, g21, g22, g23, g24, g25, g26;
	wire g27, g28, g29, g30, g31, g32, g33, g34, g35, g36, g37;
	wire g38, g39, g40, g41, g42, g43, g44, g45, g46, g47, g48;
	wire g49, g50, g51, g52, g53, g54, g55, g56, g57, g58, g59;
	wire g60, g61, g62, g63, g64, g65, g66, g67, g68, g69, g70;
	wire g71, g72, g73, g74, g75, g76, g77, g78, g79, g80, g81;
	wire g83, g84, g85, g86, g87, g88, g89, g90, g91, g92, g93;
	wire g94, g95, g96, g97, g98, g99, g100, g101, g102, g103, g104;
	wire g105, g106, g107, g108, g109, g110, g111, g112, g113, g114, g115;
	wire g116, g117, g118, g119, g120, g121, g122, g123, g124, g125, g126;
	wire g127, g128, g129, g130, g131, g683, g132, g694, g133, g134, g135;
	wire g136, g137, g138, g139, g140, g141, g142, g143, g144, g145, g146;
	wire g147, g148, g149, g150, g151, g152, g670, g153, g154, g155, g156;
	wire g157, g158, g159, g160, g161, g162, g163, g164, g165, g166, g167;
	wire g168, g169, g170, g171, g172, g173, g174, g175, g176, g177, g178;
	wire g179, g180, g181, g182, g183, g184, g185, g186, g187, g188, g189;
	wire g190, g657, g191, g192, g193, g194, g195, g196, g197, g198, g200;
	wire g201, g202, g203, g204, g205, g206, g207, g208, g209, g644, g210;
	wire g211, g212, g213, g214, g215, g216, g217, g218, g219, g220, g221;
	wire g222, g223, g224, g225, g226, g227, g228, g229, g230, g231, g232;
	wire g631, g233, g234, g235, g236, g237, g238, g239, g240, g241, g242;
	wire g243, g244, g245, g246, g247, g248, g249, g250, g251, g252, g253;
	wire g254, g255, g256, g257, g258, g259, g260, g261, g262, g264, g265;
	wire g266, g267, g268, g269, g270, g271, g272, g273, g274, g275, g276;
	wire g277, g278, g279, g280, g281, g282, g283, g284, g285, g286, g287;
	wire g288, g289, g290, g291, g292, g293, g294, g295, g296, g297, g298;
	wire g299, g300, g301, g302, g303, g304, g305, g607, g306, g307, g308;
	wire g309, g310, g311, g312, g313, g314, g315, g316, g317, g318, g319;
	wire g618, g321, g322, g596, g323, g324, g325, g326, g327, g328, g329;
	wire g330, g331, g332, g333, g334, g335, g336, g337, g338, g339, g340;
	wire g341, g342, g343, g344, g345, g346, g347, g348, g349, g350, g351;
	wire g352, g353, g354, g355, g357, g358, g359, g360, g361, g362, g363;
	wire g364, g365, g366, g367, g368, g369, g370, g371, g372, g373, g374;
	wire g375, g376, g377, g378, g379, g380, g381, g382, g383, g384, g385;
	wire g386, g387, g388, g389, g390, g391, g392, g583, g393, g394, g396;
	wire g397, g398, g399, g400, g401, g402, g403, g404, g405, g406, g407;
	wire g408, g409, g410, g411, g412, g413, g414, g415, g416, g417, g419;
	wire g420, g421, g422, g572, g423, g424, g425, g426, g427, g428, g429;
	wire g430, g431, g432, g433, g434, g435, g436, g438, g439, g440, g441;
	wire g442, g443, g444, g445, g446, g447, g448, g449, g559, g450, g451;
	wire g452, g453, g455, g456, g457, g458, g459, g460, g461, g462, g463;
	wire g464, g465, g466, g468, g469, g470, g471, g472, g473, g474, g475;
	wire g476, g477, g478, g549, g479, g480, g481, g482, g483, g484, g485;
	wire g486, g487, g488, g489, g491, g492, g493, g494, g495, g496, g497;
	wire g498, g499, g500, g501, g502, g503, g504, g505, g506, g507, g508;
	wire g509, g511, g512, g513, g514, g515, g516, g517, g543, g518, g519;
	wire g521, g522, g524, g525, g526, g527, g528, g529, g530, g531, g533;
	wire g534, g535, g536, g538, g539, g541, g544, g545, g546, g547, g548;
	wire g550, g551, g552, g554, g553, g555, g556, g557, g558, g560, g561;
	wire g562, g565, g563, g564, g568, g569, g566, g567, g570, g571, g573;
	wire g574, g575, g578, g576, g577, g580, g581, g579, g582, g584, g585;
	wire g586, g589, g587, g588, g592, g593, g590, g591, g594, g595, g597;
	wire g598, g599, g601, g600, g604, g602, g603, g605, g606, g608, g609;
	wire g610, g612, g611, g615, g613, g614, g616, g617, g619, g620, g621;
	wire g624, g622, g623, g627, g628, g625, g626, g629, g630, g632, g633;
	wire g634, g637, g635, g636, g640, g641, g638, g639, g642, g643, g645;
	wire g646, g647, g650, g648, g649, g653, g654, g651, g652, g655, g656;
	wire g658, g659, g660, g663, g661, g662, g666, g667, g664, g665, g668;
	wire g669, g671, g672, g673, g676, g674, g675, g679, g680, g677, g678;
	wire g681, g682, g684, g685, g686, g689, g687, g688, g691, g692, g690;
	wire g693, g695, g696, g697, g699, g698, g702, g700, g701, g703, g704;
	wire satCompare0, satCompare1, satCompare2, satMask0, satMask1, satCompareLevel0_0, satMaskLevel0_0, satWreckOut;


	assign g23 = (((!i_6_) & (!sk[0]) & (!i_7_) & (!i_8_)) + ((!i_6_) & (!sk[0]) & (!i_7_) & (i_8_)) + ((!i_6_) & (!sk[0]) & (i_7_) & (!i_8_)) + ((!i_6_) & (!sk[0]) & (i_7_) & (i_8_)) + ((i_6_) & (!sk[0]) & (!i_7_) & (!i_8_)) + ((i_6_) & (!sk[0]) & (!i_7_) & (i_8_)) + ((i_6_) & (!sk[0]) & (i_7_) & (i_8_)));
	assign g6 = (((i_6_) & (!sk[0]) & (!i_7_) & (i_8_)) + ((i_6_) & (sk[0]) & (!i_7_) & (!i_8_)) + ((i_6_) & (sk[0]) & (!i_7_) & (i_8_)) + ((i_6_) & (sk[0]) & (i_7_) & (!i_8_)) + ((i_6_) & (sk[0]) & (i_7_) & (i_8_)));
	assign g24 = (((!i_0_) & (!i_1_) & (!sk[1]) & (i_2_)) + ((!i_0_) & (!i_1_) & (sk[1]) & (!i_2_)) + ((!i_0_) & (!i_1_) & (sk[1]) & (i_2_)) + ((!i_0_) & (i_1_) & (!sk[1]) & (i_2_)) + ((!i_0_) & (i_1_) & (sk[1]) & (!i_2_)) + ((i_0_) & (!i_1_) & (!sk[1]) & (!i_2_)) + ((i_0_) & (!i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (!i_1_) & (sk[1]) & (!i_2_)) + ((i_0_) & (!i_1_) & (sk[1]) & (i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (!i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (i_1_) & (sk[1]) & (!i_2_)) + ((i_0_) & (i_1_) & (sk[1]) & (i_2_)));
	assign g27 = (((!i_0_) & (!i_1_) & (sk[1]) & (!i_2_)) + ((!i_0_) & (!i_1_) & (sk[1]) & (i_2_)) + ((!i_0_) & (i_1_) & (sk[1]) & (!i_2_)) + ((!i_0_) & (i_1_) & (sk[1]) & (i_2_)) + ((i_0_) & (!i_1_) & (!sk[1]) & (!i_2_)) + ((i_0_) & (!i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (!i_1_) & (sk[1]) & (!i_2_)) + ((i_0_) & (!i_1_) & (sk[1]) & (i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (!i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (i_1_) & (sk[1]) & (!i_2_)));
	assign g42 = (((!i_0_) & (!sk[1]) & (!i_1_) & (i_2_)) + ((!i_0_) & (!sk[1]) & (i_1_) & (i_2_)) + ((i_0_) & (!sk[1]) & (!i_1_) & (!i_2_)) + ((i_0_) & (!sk[1]) & (!i_1_) & (i_2_)) + ((i_0_) & (!sk[1]) & (i_1_) & (!i_2_)) + ((i_0_) & (!sk[1]) & (i_1_) & (i_2_)) + ((i_0_) & (sk[1]) & (!i_1_) & (i_2_)));
	assign g45 = (((!i_3_) & (!i_4_) & (!sk[2]) & (!i_5_)) + ((!i_3_) & (!i_4_) & (!sk[2]) & (i_5_)) + ((!i_3_) & (i_4_) & (!sk[2]) & (!i_5_)) + ((!i_3_) & (i_4_) & (!sk[2]) & (i_5_)) + ((i_3_) & (!i_4_) & (!sk[2]) & (!i_5_)) + ((i_3_) & (!i_4_) & (!sk[2]) & (i_5_)) + ((i_3_) & (i_4_) & (!sk[2]) & (i_5_)));
	assign g1 = (((!i_0_) & (!i_1_) & (!sk[1]) & (i_2_)) + ((!i_0_) & (!i_1_) & (sk[1]) & (!i_2_)) + ((!i_0_) & (!i_1_) & (sk[1]) & (i_2_)) + ((!i_0_) & (i_1_) & (!sk[1]) & (!i_2_)) + ((!i_0_) & (i_1_) & (!sk[1]) & (i_2_)) + ((!i_0_) & (i_1_) & (sk[1]) & (!i_2_)) + ((!i_0_) & (i_1_) & (sk[1]) & (i_2_)) + ((i_0_) & (!i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (!i_1_) & (sk[1]) & (i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (!i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (i_1_) & (sk[1]) & (!i_2_)) + ((i_0_) & (i_1_) & (sk[1]) & (i_2_)));
	assign g2 = (((!i_6_) & (i_7_) & (sk[0]) & (!i_8_)) + ((!i_6_) & (i_7_) & (sk[0]) & (i_8_)) + ((i_6_) & (!i_7_) & (!sk[0]) & (!i_8_)) + ((i_6_) & (i_7_) & (sk[0]) & (!i_8_)) + ((i_6_) & (i_7_) & (sk[0]) & (i_8_)));
	assign g25 = (((!i_0_) & (!i_1_) & (!sk[1]) & (i_2_)) + ((!i_0_) & (!i_1_) & (sk[1]) & (!i_2_)) + ((!i_0_) & (!i_1_) & (sk[1]) & (i_2_)) + ((!i_0_) & (i_1_) & (!sk[1]) & (!i_2_)) + ((!i_0_) & (i_1_) & (!sk[1]) & (i_2_)) + ((!i_0_) & (i_1_) & (sk[1]) & (i_2_)) + ((i_0_) & (!i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (!i_1_) & (sk[1]) & (!i_2_)) + ((i_0_) & (!i_1_) & (sk[1]) & (i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (!i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (i_1_) & (sk[1]) & (!i_2_)) + ((i_0_) & (i_1_) & (sk[1]) & (i_2_)));
	assign g21 = (((!i_3_) & (!sk[2]) & (!i_4_) & (!i_5_)) + ((!i_3_) & (!sk[2]) & (!i_4_) & (i_5_)) + ((!i_3_) & (!sk[2]) & (i_4_) & (!i_5_)) + ((!i_3_) & (!sk[2]) & (i_4_) & (i_5_)) + ((i_3_) & (!sk[2]) & (!i_4_) & (!i_5_)) + ((i_3_) & (!sk[2]) & (i_4_) & (!i_5_)) + ((i_3_) & (!sk[2]) & (i_4_) & (i_5_)));
	assign g110 = (((!i_0_) & (!i_1_) & (!sk[1]) & (i_2_)) + ((!i_0_) & (!i_1_) & (sk[1]) & (i_2_)) + ((!i_0_) & (i_1_) & (!sk[1]) & (!i_2_)) + ((!i_0_) & (i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (!i_1_) & (!sk[1]) & (i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (!i_2_)) + ((i_0_) & (i_1_) & (!sk[1]) & (i_2_)));
	assign g13 = (((!i_0_) & (!i_1_) & (sk[3]) & (!i_2_)) + ((!i_0_) & (!i_1_) & (sk[3]) & (i_2_)) + ((!i_0_) & (i_1_) & (!sk[3]) & (!i_2_)) + ((!i_0_) & (i_1_) & (!sk[3]) & (i_2_)) + ((!i_0_) & (i_1_) & (sk[3]) & (!i_2_)) + ((!i_0_) & (i_1_) & (sk[3]) & (i_2_)) + ((i_0_) & (!i_1_) & (!sk[3]) & (!i_2_)) + ((i_0_) & (!i_1_) & (!sk[3]) & (i_2_)) + ((i_0_) & (!i_1_) & (sk[3]) & (!i_2_)) + ((i_0_) & (!i_1_) & (sk[3]) & (i_2_)) + ((i_0_) & (i_1_) & (!sk[3]) & (!i_2_)) + ((i_0_) & (i_1_) & (!sk[3]) & (i_2_)) + ((i_0_) & (i_1_) & (sk[3]) & (i_2_)));
	assign g28 = (((!sk[0]) & (i_6_) & (i_7_) & (i_8_)) + ((sk[0]) & (!i_6_) & (!i_7_) & (i_8_)) + ((sk[0]) & (!i_6_) & (i_7_) & (i_8_)) + ((sk[0]) & (i_6_) & (!i_7_) & (!i_8_)) + ((sk[0]) & (i_6_) & (!i_7_) & (i_8_)) + ((sk[0]) & (i_6_) & (i_7_) & (!i_8_)) + ((sk[0]) & (i_6_) & (i_7_) & (i_8_)));
	assign g12 = (((!i_6_) & (!sk[0]) & (i_7_) & (!i_8_)) + ((!i_6_) & (sk[0]) & (!i_7_) & (i_8_)) + ((!i_6_) & (sk[0]) & (i_7_) & (i_8_)) + ((i_6_) & (sk[0]) & (!i_7_) & (i_8_)) + ((i_6_) & (sk[0]) & (i_7_) & (i_8_)));
	assign g11 = (((!sk[2]) & (!i_3_) & (!i_4_) & (!i_5_)) + ((!sk[2]) & (!i_3_) & (i_4_) & (!i_5_)) + ((!sk[2]) & (!i_3_) & (i_4_) & (i_5_)) + ((!sk[2]) & (i_3_) & (!i_4_) & (!i_5_)) + ((!sk[2]) & (i_3_) & (!i_4_) & (i_5_)) + ((!sk[2]) & (i_3_) & (i_4_) & (!i_5_)) + ((!sk[2]) & (i_3_) & (i_4_) & (i_5_)));
	assign g35 = (((!i_6_) & (!sk[0]) & (!i_7_) & (!i_8_)));
	assign g36 = (((!i_3_) & (!i_4_) & (!sk[2]) & (!i_5_)) + ((!i_3_) & (!i_4_) & (!sk[2]) & (i_5_)) + ((!i_3_) & (i_4_) & (!sk[2]) & (!i_5_)) + ((!i_3_) & (i_4_) & (!sk[2]) & (i_5_)) + ((i_3_) & (!i_4_) & (!sk[2]) & (i_5_)) + ((i_3_) & (i_4_) & (!sk[2]) & (!i_5_)) + ((i_3_) & (i_4_) & (!sk[2]) & (i_5_)));
	assign g38 = (((!sk[2]) & (!i_3_) & (!i_4_) & (!i_5_)) + ((!sk[2]) & (!i_3_) & (!i_4_) & (i_5_)) + ((!sk[2]) & (!i_3_) & (i_4_) & (!i_5_)) + ((!sk[2]) & (i_3_) & (!i_4_) & (!i_5_)) + ((!sk[2]) & (i_3_) & (!i_4_) & (i_5_)) + ((!sk[2]) & (i_3_) & (i_4_) & (!i_5_)) + ((!sk[2]) & (i_3_) & (i_4_) & (i_5_)));
	assign g8 = (((!i_6_) & (i_7_) & (!sk[3]) & (!i_8_)) + ((!i_6_) & (i_7_) & (!sk[3]) & (i_8_)) + ((!i_6_) & (i_7_) & (sk[3]) & (i_8_)) + ((i_6_) & (!i_7_) & (!sk[3]) & (!i_8_)) + ((i_6_) & (!i_7_) & (!sk[3]) & (i_8_)) + ((i_6_) & (i_7_) & (!sk[3]) & (!i_8_)) + ((i_6_) & (i_7_) & (!sk[3]) & (i_8_)));
	assign g32 = (((!sk[2]) & (!i_3_) & (!i_4_) & (!i_5_)));
	assign g3 = (((!i_3_) & (!sk[3]) & (i_4_) & (!i_5_)) + ((!i_3_) & (!sk[3]) & (i_4_) & (i_5_)) + ((!i_3_) & (sk[3]) & (i_4_) & (!i_5_)) + ((i_3_) & (!sk[3]) & (!i_4_) & (!i_5_)) + ((i_3_) & (!sk[3]) & (!i_4_) & (i_5_)) + ((i_3_) & (!sk[3]) & (i_4_) & (!i_5_)) + ((i_3_) & (!sk[3]) & (i_4_) & (i_5_)));
	assign g48 = (((!i_6_) & (!sk[3]) & (g47)) + ((!i_6_) & (sk[3]) & (g47)) + ((i_6_) & (!sk[3]) & (g47)));
	assign g59 = (((!i_3_) & (!sk[4]) & (!i_4_) & (!i_5_)) + ((!i_3_) & (!sk[4]) & (!i_4_) & (i_5_)) + ((!i_3_) & (!sk[4]) & (i_4_) & (!i_5_)) + ((!i_3_) & (!sk[4]) & (i_4_) & (i_5_)) + ((i_3_) & (!sk[4]) & (!i_4_) & (!i_5_)) + ((i_3_) & (!sk[4]) & (!i_4_) & (i_5_)) + ((i_3_) & (!sk[4]) & (i_4_) & (!i_5_)));
	assign g47 = (((!i_7_) & (!sk[5]) & (i_8_)) + ((!i_7_) & (sk[5]) & (i_8_)) + ((i_7_) & (sk[5]) & (i_8_)));
	assign g63 = (((!i_7_) & (!sk[5]) & (!i_8_)));
	assign g50 = (((!sk[4]) & (!i_4_) & (i_5_)) + ((sk[4]) & (i_4_) & (!i_5_)) + ((sk[4]) & (i_4_) & (i_5_)));
	assign g14 = (((i_7_) & (!sk[5]) & (i_8_)) + ((i_7_) & (sk[5]) & (!i_8_)) + ((i_7_) & (sk[5]) & (i_8_)));
	assign g121 = (((!sk[6]) & (!g28) & (g13)) + ((!sk[6]) & (g28) & (g13)) + ((sk[6]) & (g28) & (!g13)));
	assign g26 = (((!sk[6]) & (g11) & (g25)) + ((sk[6]) & (!g11) & (!g25)));
	assign g29 = (((g28) & (!sk[6]) & (!g1)) + ((g28) & (!sk[6]) & (g1)) + ((g28) & (sk[6]) & (!g1)));
	assign g75 = (((!g24) & (sk[6]) & (!g59)) + ((g24) & (!sk[6]) & (!g59)) + ((g24) & (!sk[6]) & (g59)));
	assign g137 = (((!sk[5]) & (i_7_) & (!i_8_)) + ((sk[5]) & (i_7_) & (!i_8_)) + ((sk[5]) & (i_7_) & (i_8_)));
	assign g184 = (((!sk[7]) & (!g59) & (g110)) + ((sk[7]) & (g59) & (!g110)) + ((sk[7]) & (g59) & (g110)));
	assign g64 = (((!i_4_) & (!i_5_) & (sk[4]) & (i_6_)) + ((!i_4_) & (i_5_) & (sk[4]) & (i_6_)) + ((i_4_) & (!i_5_) & (!sk[4]) & (!i_6_)) + ((i_4_) & (!i_5_) & (sk[4]) & (i_6_)) + ((i_4_) & (i_5_) & (sk[4]) & (i_6_)));
	assign g105 = (((!sk[8]) & (!g24) & (g38)) + ((!sk[8]) & (g24) & (!g38)) + ((!sk[8]) & (g24) & (g38)) + ((sk[8]) & (g24) & (!g38)) + ((sk[8]) & (g24) & (g38)));
	assign g189 = (((!sk[7]) & (g3) & (g110)) + ((sk[7]) & (g3) & (!g110)) + ((sk[7]) & (g3) & (g110)));
	assign g4 = (((!sk[9]) & (g2) & (g3)) + ((sk[9]) & (!g2) & (g3)) + ((sk[9]) & (g2) & (g3)));
	assign g5 = (((!i_3_) & (!sk[4]) & (i_4_)) + ((i_3_) & (sk[4]) & (!i_4_)) + ((i_3_) & (sk[4]) & (i_4_)));
	assign g46 = (((!g25) & (!sk[9]) & (!g45)));
	assign g77 = (((!sk[7]) & (!g25) & (!g59)));
	assign g99 = (((!sk[9]) & (!g25) & (g3)) + ((sk[9]) & (!g25) & (g3)) + ((sk[9]) & (g25) & (g3)));
	assign g127 = (((!i_0_) & (!sk[3]) & (i_1_)) + ((i_0_) & (!sk[3]) & (i_1_)) + ((i_0_) & (sk[3]) & (i_1_)));
	assign g129 = (((!sk[9]) & (g42) & (g32)) + ((sk[9]) & (!g42) & (g32)) + ((sk[9]) & (g42) & (g32)));
	assign g243 = (((!g25) & (!sk[9]) & (!g36)));
	assign g7 = (((!g1) & (!sk[10]) & (g6)) + ((g1) & (sk[10]) & (!g6)) + ((g1) & (sk[10]) & (g6)));
	assign g41 = (((!g27) & (!sk[10]) & (g35)) + ((!g27) & (sk[10]) & (g35)) + ((g27) & (sk[10]) & (g35)));
	assign g161 = (((!g11) & (!sk[7]) & (g110)) + ((g11) & (sk[7]) & (!g110)) + ((g11) & (sk[7]) & (g110)));
	assign g181 = (((!sk[7]) & (!g45) & (g110)) + ((sk[7]) & (g45) & (!g110)) + ((sk[7]) & (g45) & (g110)));
	assign g194 = (((!sk[10]) & (!g21) & (g6)) + ((sk[10]) & (g21) & (!g6)) + ((sk[10]) & (g21) & (g6)));
	assign g22 = (((!sk[9]) & (!g21) & (g2)) + ((sk[9]) & (g21) & (!g2)) + ((sk[9]) & (g21) & (g2)));
	assign g33 = (((!g24) & (!sk[8]) & (g3)) + ((g24) & (sk[8]) & (g3)));
	assign g37 = (((!i_6_) & (!sk[5]) & (!i_7_)));
	assign g60 = (((i_6_) & (!sk[5]) & (i_7_)) + ((i_6_) & (sk[5]) & (i_7_)));
	assign g70 = (((!sk[10]) & (!g25) & (g32)) + ((sk[10]) & (!g25) & (g32)) + ((sk[10]) & (g25) & (g32)));
	assign g88 = (((!g42) & (sk[10]) & (g36)) + ((g42) & (!sk[10]) & (!g36)) + ((g42) & (sk[10]) & (g36)));
	assign g98 = (((!sk[8]) & (!g24) & (!g36)));
	assign g49 = (((!g32) & (!sk[6]) & (g13)) + ((g32) & (!sk[6]) & (g13)) + ((g32) & (sk[6]) & (!g13)));
	assign g71 = (((!g42) & (sk[7]) & (g59)) + ((g42) & (!sk[7]) & (!g59)) + ((g42) & (sk[7]) & (g59)));
	assign g141 = (((!sk[8]) & (g35) & (!g24)) + ((sk[8]) & (g35) & (!g24)) + ((sk[8]) & (g35) & (g24)));
	assign g9 = (((!sk[10]) & (g8) & (!g1)) + ((sk[10]) & (g8) & (!g1)) + ((sk[10]) & (g8) & (g1)));
	assign g73 = (((!sk[8]) & (!g11) & (!g24)));
	assign g84 = (((!sk[8]) & (!g1) & (!g38)));
	assign g85 = (((!i_4_) & (!i_5_) & (!sk[4]) & (i_6_)) + ((!i_4_) & (!i_5_) & (sk[4]) & (i_6_)) + ((!i_4_) & (i_5_) & (sk[4]) & (i_6_)) + ((i_4_) & (!i_5_) & (sk[4]) & (i_6_)) + ((i_4_) & (i_5_) & (sk[4]) & (i_6_)));
	assign g91 = (((!sk[6]) & (g36) & (!g13)) + ((!sk[6]) & (g36) & (g13)) + ((sk[6]) & (!g36) & (!g13)));
	assign g111 = (((!sk[11]) & (i_6_) & (!i_7_)) + ((!sk[11]) & (i_6_) & (i_7_)) + ((sk[11]) & (!i_6_) & (i_7_)));
	assign g116 = (((i_3_) & (!sk[4]) & (i_5_)) + ((i_3_) & (sk[4]) & (!i_5_)) + ((i_3_) & (sk[4]) & (i_5_)));
	assign g123 = (((g50) & (!sk[11]) & (!g8)) + ((g50) & (!sk[11]) & (g8)) + ((g50) & (sk[11]) & (g8)));
	assign g134 = (((!i_4_) & (!sk[11]) & (!i_5_) & (i_6_)) + ((!i_4_) & (!sk[11]) & (i_5_) & (!i_6_)) + ((!i_4_) & (!sk[11]) & (i_5_) & (i_6_)) + ((!i_4_) & (sk[11]) & (!i_5_) & (!i_6_)) + ((i_4_) & (!sk[11]) & (!i_5_) & (i_6_)) + ((i_4_) & (!sk[11]) & (i_5_) & (!i_6_)) + ((i_4_) & (!sk[11]) & (i_5_) & (i_6_)));
	assign g159 = (((!g21) & (sk[11]) & (g48)) + ((g21) & (!sk[11]) & (g48)));
	assign g265 = (((!sk[11]) & (!g27) & (!i_6_) & (g47)) + ((!sk[11]) & (!g27) & (i_6_) & (g47)) + ((!sk[11]) & (g27) & (!i_6_) & (g47)) + ((!sk[11]) & (g27) & (i_6_) & (g47)) + ((sk[11]) & (!g27) & (!i_6_) & (g47)));
	assign g359 = (((!sk[11]) & (g21) & (!g110)) + ((!sk[11]) & (g21) & (g110)) + ((sk[11]) & (!g21) & (g110)));
	assign g472 = (((!sk[3]) & (!i_3_) & (!i_0_) & (i_1_)) + ((!sk[3]) & (!i_3_) & (i_0_) & (!i_1_)) + ((!sk[3]) & (!i_3_) & (i_0_) & (i_1_)) + ((!sk[3]) & (i_3_) & (!i_0_) & (i_1_)) + ((!sk[3]) & (i_3_) & (i_0_) & (!i_1_)) + ((!sk[3]) & (i_3_) & (i_0_) & (i_1_)) + ((sk[3]) & (!i_3_) & (!i_0_) & (!i_1_)));
	assign g15 = (((i_4_) & (i_5_) & (!i_6_)));
	assign g16 = (((g14) & (g15)));
	assign g51 = (((!i_3_) & (i_0_) & (!i_2_)));
	assign g67 = (((!g27) & (g2)));
	assign g117 = (((!g13) & (g116)));
	assign g230 = (((!i_3_) & (i_1_) & (i_2_)));
	assign g94 = (((!i_3_) & (i_0_) & (!i_1_)));
	assign g100 = (((g3) & (!g13)));
	assign g135 = (((i_3_) & (i_2_) & (g47) & (g134)));
	assign g158 = (((!g1) & (!g59)));
	assign g219 = (((g63) & (g15)));
	assign g392 = (((!i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (!g8) & (!g117)) + ((!i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (!g8) & (g117)) + ((!i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (g8) & (!g117)) + ((!i_4_) & (!i_5_) & (!i_0_) & (i_1_) & (!g8) & (!g117)) + ((!i_4_) & (!i_5_) & (!i_0_) & (i_1_) & (!g8) & (g117)) + ((!i_4_) & (!i_5_) & (i_0_) & (!i_1_) & (!g8) & (!g117)) + ((!i_4_) & (!i_5_) & (i_0_) & (!i_1_) & (!g8) & (g117)) + ((!i_4_) & (!i_5_) & (i_0_) & (!i_1_) & (g8) & (!g117)) + ((!i_4_) & (!i_5_) & (i_0_) & (i_1_) & (!g8) & (!g117)) + ((!i_4_) & (!i_5_) & (i_0_) & (i_1_) & (!g8) & (g117)) + ((!i_4_) & (i_5_) & (!i_0_) & (!i_1_) & (!g8) & (!g117)) + ((!i_4_) & (i_5_) & (!i_0_) & (!i_1_) & (!g8) & (g117)) + ((!i_4_) & (i_5_) & (!i_0_) & (!i_1_) & (g8) & (!g117)) + ((!i_4_) & (i_5_) & (!i_0_) & (i_1_) & (!g8) & (!g117)) + ((!i_4_) & (i_5_) & (!i_0_) & (i_1_) & (!g8) & (g117)) + ((!i_4_) & (i_5_) & (!i_0_) & (i_1_) & (g8) & (!g117)) + ((!i_4_) & (i_5_) & (i_0_) & (!i_1_) & (!g8) & (!g117)) + ((!i_4_) & (i_5_) & (i_0_) & (!i_1_) & (!g8) & (g117)) + ((!i_4_) & (i_5_) & (i_0_) & (i_1_) & (!g8) & (!g117)) + ((!i_4_) & (i_5_) & (i_0_) & (i_1_) & (!g8) & (g117)) + ((!i_4_) & (i_5_) & (i_0_) & (i_1_) & (g8) & (!g117)) + ((i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (!g8) & (!g117)) + ((i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (!g8) & (g117)) + ((i_4_) & (!i_5_) & (!i_0_) & (!i_1_) & (g8) & (!g117)) + ((i_4_) & (!i_5_) & (!i_0_) & (i_1_) & (!g8) & (!g117)) + ((i_4_) & (!i_5_) & (!i_0_) & (i_1_) & (!g8) & (g117)) + ((i_4_) & (!i_5_) & (!i_0_) & (i_1_) & (g8) & (!g117)) + ((i_4_) & (!i_5_) & (i_0_) & (!i_1_) & (!g8) & (!g117)) + ((i_4_) & (!i_5_) & (i_0_) & (!i_1_) & (!g8) & (g117)) + ((i_4_) & (!i_5_) & (i_0_) & (!i_1_) & (g8) & (!g117)) + ((i_4_) & (!i_5_) & (i_0_) & (i_1_) & (!g8) & (!g117)) + ((i_4_) & (!i_5_) & (i_0_) & (i_1_) & (!g8) & (g117)) + ((i_4_) & (!i_5_) & (i_0_) & (i_1_) & (g8) & (!g117)) + ((i_4_) & (i_5_) & (!i_0_) & (!i_1_) & (!g8) & (!g117)) + ((i_4_) & (i_5_) & (!i_0_) & (!i_1_) & (!g8) & (g117)) + ((i_4_) & (i_5_) & (!i_0_) & (!i_1_) & (g8) & (!g117)) + ((i_4_) & (i_5_) & (!i_0_) & (i_1_) & (!g8) & (!g117)) + ((i_4_) & (i_5_) & (!i_0_) & (i_1_) & (!g8) & (g117)) + ((i_4_) & (i_5_) & (!i_0_) & (i_1_) & (g8) & (!g117)) + ((i_4_) & (i_5_) & (i_0_) & (!i_1_) & (!g8) & (!g117)) + ((i_4_) & (i_5_) & (i_0_) & (!i_1_) & (!g8) & (g117)) + ((i_4_) & (i_5_) & (i_0_) & (!i_1_) & (g8) & (!g117)) + ((i_4_) & (i_5_) & (i_0_) & (i_1_) & (!g8) & (!g117)) + ((i_4_) & (i_5_) & (i_0_) & (i_1_) & (!g8) & (g117)) + ((i_4_) & (i_5_) & (i_0_) & (i_1_) & (g8) & (!g117)));
	assign g447 = (((!g14) & (!g24) & (!g64) & (!g194) & (!g446)) + ((!g14) & (!g24) & (g64) & (!g194) & (!g446)) + ((!g14) & (g24) & (!g64) & (!g194) & (!g446)) + ((!g14) & (g24) & (!g64) & (g194) & (!g446)) + ((!g14) & (g24) & (g64) & (!g194) & (!g446)) + ((!g14) & (g24) & (g64) & (g194) & (!g446)) + ((g14) & (!g24) & (!g64) & (!g194) & (!g446)) + ((g14) & (g24) & (!g64) & (!g194) & (!g446)) + ((g14) & (g24) & (!g64) & (g194) & (!g446)) + ((g14) & (g24) & (g64) & (!g194) & (!g446)) + ((g14) & (g24) & (g64) & (g194) & (!g446)));
	assign g448 = (((!g25) & (!g2) & (!g38) & (!g110)) + ((!g25) & (!g2) & (!g38) & (g110)) + ((!g25) & (!g2) & (g38) & (!g110)) + ((!g25) & (!g2) & (g38) & (g110)) + ((!g25) & (g2) & (g38) & (!g110)) + ((!g25) & (g2) & (g38) & (g110)) + ((g25) & (!g2) & (!g38) & (!g110)) + ((g25) & (!g2) & (!g38) & (g110)) + ((g25) & (!g2) & (g38) & (!g110)) + ((g25) & (!g2) & (g38) & (g110)) + ((g25) & (g2) & (!g38) & (!g110)) + ((g25) & (g2) & (g38) & (!g110)) + ((g25) & (g2) & (g38) & (g110)));
	assign g449 = (((!i_5_) & (!g6) & (!g23) & (!g110) & (!g440)) + ((!i_5_) & (!g6) & (!g23) & (g110) & (!g440)) + ((!i_5_) & (!g6) & (g23) & (!g110) & (!g440)) + ((!i_5_) & (!g6) & (g23) & (!g110) & (g440)) + ((!i_5_) & (!g6) & (g23) & (g110) & (!g440)) + ((!i_5_) & (!g6) & (g23) & (g110) & (g440)) + ((!i_5_) & (g6) & (!g23) & (!g110) & (!g440)) + ((!i_5_) & (g6) & (g23) & (!g110) & (!g440)) + ((!i_5_) & (g6) & (g23) & (!g110) & (g440)) + ((i_5_) & (!g6) & (!g23) & (!g110) & (!g440)) + ((i_5_) & (!g6) & (!g23) & (!g110) & (g440)) + ((i_5_) & (!g6) & (!g23) & (g110) & (!g440)) + ((i_5_) & (!g6) & (!g23) & (g110) & (g440)) + ((i_5_) & (!g6) & (g23) & (!g110) & (!g440)) + ((i_5_) & (!g6) & (g23) & (!g110) & (g440)) + ((i_5_) & (!g6) & (g23) & (g110) & (!g440)) + ((i_5_) & (!g6) & (g23) & (g110) & (g440)) + ((i_5_) & (g6) & (!g23) & (!g110) & (!g440)) + ((i_5_) & (g6) & (!g23) & (!g110) & (g440)) + ((i_5_) & (g6) & (!g23) & (g110) & (!g440)) + ((i_5_) & (g6) & (!g23) & (g110) & (g440)) + ((i_5_) & (g6) & (g23) & (!g110) & (!g440)) + ((i_5_) & (g6) & (g23) & (!g110) & (g440)) + ((i_5_) & (g6) & (g23) & (g110) & (!g440)) + ((i_5_) & (g6) & (g23) & (g110) & (g440)));
	assign g17 = (((i_3_) & (i_0_) & (!i_2_)));
	assign g18 = (((g16) & (g17)));
	assign g43 = (((!g21) & (g28) & (g42)));
	assign g57 = (((i_3_) & (!i_1_) & (i_2_)));
	assign g65 = (((i_3_) & (i_0_) & (!i_1_) & (g64)));
	assign g86 = (((i_3_) & (i_0_) & (i_2_)));
	assign g90 = (((!g45) & (!g6) & (!g13) & (!g89)) + ((!g45) & (!g6) & (g13) & (!g89)) + ((!g45) & (g6) & (g13) & (!g89)) + ((g45) & (!g6) & (!g13) & (!g89)) + ((g45) & (!g6) & (g13) & (!g89)) + ((g45) & (g6) & (!g13) & (!g89)) + ((g45) & (g6) & (g13) & (!g89)));
	assign g95 = (((g47) & (g94)));
	assign g120 = (((i_3_) & (i_4_)));
	assign g150 = (((g12) & (!g59) & (!g13)));
	assign g155 = (((!g11) & (!g27) & (g28)));
	assign g167 = (((g14) & (g134)));
	assign g212 = (((!g45) & (!g23) & (!g24)));
	assign g217 = (((!i_3_) & (i_5_) & (!i_6_)));
	assign g225 = (((!i_3_) & (!i_4_) & (!i_6_)));
	assign g252 = (((!g27) & (g28) & (!g45)));
	assign g290 = (((g42) & (g2) & (!g38)));
	assign g294 = (((g28) & (!g45) & (!g24)));
	assign g296 = (((g8) & (g243)));
	assign g401 = (((!i_3_) & (g50) & (!i_0_) & (i_2_) & (!i_6_)));
	assign g440 = (((!i_3_) & (!i_1_) & (i_2_)));
	assign g20 = (((!g1) & (!g4) & (!g10) & (g19)) + ((g1) & (!g4) & (!g10) & (g19)) + ((g1) & (g4) & (!g10) & (g19)));
	assign g30 = (((!g11) & (!g27) & (!g21) & (!g6) & (g29)) + ((!g11) & (!g27) & (!g21) & (g6) & (!g29)) + ((!g11) & (!g27) & (!g21) & (g6) & (g29)) + ((!g11) & (!g27) & (g21) & (g6) & (!g29)) + ((!g11) & (!g27) & (g21) & (g6) & (g29)) + ((!g11) & (g27) & (!g21) & (!g6) & (g29)) + ((!g11) & (g27) & (!g21) & (g6) & (g29)) + ((g11) & (!g27) & (!g21) & (!g6) & (g29)) + ((g11) & (!g27) & (!g21) & (g6) & (g29)) + ((g11) & (g27) & (!g21) & (!g6) & (g29)) + ((g11) & (g27) & (!g21) & (g6) & (g29)));
	assign g31 = (((!g22) & (!g23) & (!g24) & (!g26) & (!g30)) + ((!g22) & (!g23) & (g24) & (!g26) & (!g30)) + ((!g22) & (g23) & (!g24) & (!g26) & (!g30)) + ((!g22) & (g23) & (!g24) & (g26) & (!g30)) + ((!g22) & (g23) & (g24) & (!g26) & (!g30)) + ((!g22) & (g23) & (g24) & (g26) & (!g30)) + ((g22) & (!g23) & (g24) & (!g26) & (!g30)) + ((g22) & (g23) & (g24) & (!g26) & (!g30)) + ((g22) & (g23) & (g24) & (g26) & (!g30)));
	assign g34 = (((!g11) & (!g27) & (!g6) & (!g23) & (!g32) & (!g33)) + ((!g11) & (!g27) & (!g6) & (!g23) & (!g32) & (g33)) + ((!g11) & (!g27) & (!g6) & (!g23) & (g32) & (!g33)) + ((!g11) & (!g27) & (!g6) & (!g23) & (g32) & (g33)) + ((!g11) & (!g27) & (g6) & (!g23) & (!g32) & (!g33)) + ((!g11) & (!g27) & (g6) & (!g23) & (!g32) & (g33)) + ((!g11) & (!g27) & (g6) & (!g23) & (g32) & (!g33)) + ((!g11) & (!g27) & (g6) & (!g23) & (g32) & (g33)) + ((!g11) & (!g27) & (g6) & (g23) & (g32) & (!g33)) + ((!g11) & (!g27) & (g6) & (g23) & (g32) & (g33)) + ((!g11) & (g27) & (!g6) & (!g23) & (!g32) & (g33)) + ((!g11) & (g27) & (!g6) & (!g23) & (g32) & (g33)) + ((!g11) & (g27) & (g6) & (!g23) & (!g32) & (g33)) + ((!g11) & (g27) & (g6) & (!g23) & (g32) & (g33)) + ((g11) & (!g27) & (!g6) & (!g23) & (!g32) & (g33)) + ((g11) & (!g27) & (!g6) & (!g23) & (g32) & (g33)) + ((g11) & (!g27) & (g6) & (!g23) & (!g32) & (g33)) + ((g11) & (!g27) & (g6) & (!g23) & (g32) & (!g33)) + ((g11) & (!g27) & (g6) & (!g23) & (g32) & (g33)) + ((g11) & (!g27) & (g6) & (g23) & (g32) & (!g33)) + ((g11) & (!g27) & (g6) & (g23) & (g32) & (g33)) + ((g11) & (g27) & (!g6) & (!g23) & (!g32) & (g33)) + ((g11) & (g27) & (!g6) & (!g23) & (g32) & (g33)) + ((g11) & (g27) & (g6) & (!g23) & (!g32) & (g33)) + ((g11) & (g27) & (g6) & (!g23) & (g32) & (g33)));
	assign g40 = (((!g35) & (!g1) & (!g36) & (!g39)) + ((!g35) & (!g1) & (g36) & (!g39)) + ((!g35) & (g1) & (!g36) & (!g39)) + ((!g35) & (g1) & (g36) & (!g39)) + ((g35) & (!g1) & (g36) & (!g39)) + ((g35) & (g1) & (!g36) & (!g39)) + ((g35) & (g1) & (g36) & (!g39)));
	assign g52 = (((g50) & (g51)));
	assign g66 = (((!g42) & (!g45) & (!g23) & (!g36) & (g29)) + ((!g42) & (!g45) & (g23) & (!g36) & (g29)) + ((!g42) & (g45) & (!g23) & (!g36) & (g29)) + ((!g42) & (g45) & (g23) & (!g36) & (g29)) + ((g42) & (!g45) & (!g23) & (!g36) & (!g29)) + ((g42) & (!g45) & (!g23) & (!g36) & (g29)) + ((g42) & (!g45) & (!g23) & (g36) & (!g29)) + ((g42) & (!g45) & (!g23) & (g36) & (g29)) + ((g42) & (!g45) & (g23) & (!g36) & (g29)) + ((g42) & (g45) & (!g23) & (!g36) & (g29)) + ((g42) & (g45) & (g23) & (!g36) & (g29)));
	assign g69 = (((!g42) & (!g45) & (!g6) & (!g68)) + ((!g42) & (!g45) & (g6) & (!g68)) + ((!g42) & (g45) & (!g6) & (!g68)) + ((!g42) & (g45) & (g6) & (!g68)) + ((g42) & (!g45) & (!g6) & (!g68)) + ((g42) & (g45) & (!g6) & (!g68)) + ((g42) & (g45) & (g6) & (!g68)));
	assign g72 = (((!g27) & (!g28) & (!g32) & (g37) & (g71)) + ((!g27) & (!g28) & (g32) & (g37) & (g71)) + ((!g27) & (g28) & (!g32) & (g37) & (g71)) + ((!g27) & (g28) & (g32) & (!g37) & (!g71)) + ((!g27) & (g28) & (g32) & (!g37) & (g71)) + ((!g27) & (g28) & (g32) & (g37) & (!g71)) + ((!g27) & (g28) & (g32) & (g37) & (g71)) + ((g27) & (!g28) & (!g32) & (g37) & (g71)) + ((g27) & (!g28) & (g32) & (g37) & (g71)) + ((g27) & (g28) & (!g32) & (g37) & (g71)) + ((g27) & (g28) & (g32) & (g37) & (g71)));
	assign g74 = (((g6) & (!g24) & (g32)));
	assign g80 = (((!g21) & (!g8) & (!g24) & (g69) & (g79)) + ((!g21) & (!g8) & (g24) & (g69) & (g79)) + ((!g21) & (g8) & (g24) & (g69) & (g79)) + ((g21) & (!g8) & (!g24) & (g69) & (g79)) + ((g21) & (!g8) & (g24) & (g69) & (g79)) + ((g21) & (g8) & (!g24) & (g69) & (g79)) + ((g21) & (g8) & (g24) & (g69) & (g79)));
	assign g83 = (((!g21) & (!g8) & (!g24) & (!g77) & (g37)) + ((!g21) & (!g8) & (!g24) & (g77) & (g37)) + ((!g21) & (g8) & (!g24) & (!g77) & (g37)) + ((!g21) & (g8) & (!g24) & (g77) & (!g37)) + ((!g21) & (g8) & (!g24) & (g77) & (g37)) + ((!g21) & (g8) & (g24) & (g77) & (!g37)) + ((!g21) & (g8) & (g24) & (g77) & (g37)) + ((g21) & (g8) & (!g24) & (g77) & (!g37)) + ((g21) & (g8) & (!g24) & (g77) & (g37)) + ((g21) & (g8) & (g24) & (g77) & (!g37)) + ((g21) & (g8) & (g24) & (g77) & (g37)));
	assign g87 = (((!g63) & (g8) & (g84) & (!g85) & (!g86)) + ((!g63) & (g8) & (g84) & (!g85) & (g86)) + ((!g63) & (g8) & (g84) & (g85) & (!g86)) + ((!g63) & (g8) & (g84) & (g85) & (g86)) + ((g63) & (!g8) & (!g84) & (g85) & (g86)) + ((g63) & (!g8) & (g84) & (g85) & (g86)) + ((g63) & (g8) & (!g84) & (g85) & (g86)) + ((g63) & (g8) & (g84) & (!g85) & (!g86)) + ((g63) & (g8) & (g84) & (!g85) & (g86)) + ((g63) & (g8) & (g84) & (g85) & (!g86)) + ((g63) & (g8) & (g84) & (g85) & (g86)));
	assign g92 = (((g42) & (g12) & (g3)));
	assign g93 = (((!g41) & (!g45) & (!g48) & (!g91) & (!g92)) + ((!g41) & (!g45) & (!g48) & (g91) & (!g92)) + ((!g41) & (!g45) & (g48) & (!g91) & (!g92)) + ((!g41) & (g45) & (!g48) & (!g91) & (!g92)) + ((!g41) & (g45) & (!g48) & (g91) & (!g92)) + ((!g41) & (g45) & (g48) & (!g91) & (!g92)) + ((g41) & (g45) & (!g48) & (!g91) & (!g92)) + ((g41) & (g45) & (!g48) & (g91) & (!g92)) + ((g41) & (g45) & (g48) & (!g91) & (!g92)));
	assign g96 = (((g85) & (g95)));
	assign g97 = (((!g27) & (!g23) & (g32)));
	assign g101 = (((!i_6_) & (!i_7_) & (i_8_) & (!g98) & (g99) & (!g100)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g98) & (g99) & (g100)) + ((!i_6_) & (!i_7_) & (i_8_) & (g98) & (g99) & (!g100)) + ((!i_6_) & (!i_7_) & (i_8_) & (g98) & (g99) & (g100)) + ((!i_6_) & (i_7_) & (!i_8_) & (g98) & (!g99) & (!g100)) + ((!i_6_) & (i_7_) & (!i_8_) & (g98) & (!g99) & (g100)) + ((!i_6_) & (i_7_) & (!i_8_) & (g98) & (g99) & (!g100)) + ((!i_6_) & (i_7_) & (!i_8_) & (g98) & (g99) & (g100)) + ((!i_6_) & (i_7_) & (i_8_) & (g98) & (!g99) & (!g100)) + ((!i_6_) & (i_7_) & (i_8_) & (g98) & (!g99) & (g100)) + ((!i_6_) & (i_7_) & (i_8_) & (g98) & (g99) & (!g100)) + ((!i_6_) & (i_7_) & (i_8_) & (g98) & (g99) & (g100)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g98) & (!g99) & (g100)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g98) & (g99) & (g100)) + ((i_6_) & (!i_7_) & (!i_8_) & (g98) & (!g99) & (g100)) + ((i_6_) & (!i_7_) & (!i_8_) & (g98) & (g99) & (g100)) + ((i_6_) & (!i_7_) & (i_8_) & (!g98) & (!g99) & (g100)) + ((i_6_) & (!i_7_) & (i_8_) & (!g98) & (g99) & (g100)) + ((i_6_) & (!i_7_) & (i_8_) & (g98) & (!g99) & (g100)) + ((i_6_) & (!i_7_) & (i_8_) & (g98) & (g99) & (g100)));
	assign g102 = (((!g8) & (g12) & (!g75) & (g49)) + ((!g8) & (g12) & (g75) & (g49)) + ((g8) & (!g12) & (g75) & (!g49)) + ((g8) & (!g12) & (g75) & (g49)) + ((g8) & (g12) & (!g75) & (g49)) + ((g8) & (g12) & (g75) & (!g49)) + ((g8) & (g12) & (g75) & (g49)));
	assign g109 = (((!g83) & (!g87) & (g90) & (g93) & (g108)));
	assign g119 = (((!g28) & (!g48) & (!g26) & (!g117) & (!g118)) + ((!g28) & (!g48) & (!g26) & (g117) & (!g118)) + ((!g28) & (!g48) & (g26) & (!g117) & (!g118)) + ((!g28) & (!g48) & (g26) & (g117) & (!g118)) + ((!g28) & (g48) & (!g26) & (!g117) & (!g118)) + ((!g28) & (g48) & (g26) & (!g117) & (!g118)) + ((g28) & (!g48) & (!g26) & (!g117) & (!g118)) + ((g28) & (!g48) & (!g26) & (g117) & (!g118)) + ((g28) & (g48) & (!g26) & (!g117) & (!g118)));
	assign g122 = (((!g42) & (!g45) & (!g6) & (!g24) & (!g3) & (g111)) + ((!g42) & (!g45) & (!g6) & (!g24) & (g3) & (g111)) + ((!g42) & (!g45) & (g6) & (!g24) & (!g3) & (g111)) + ((!g42) & (!g45) & (g6) & (!g24) & (g3) & (g111)) + ((g42) & (!g45) & (!g6) & (!g24) & (!g3) & (g111)) + ((g42) & (!g45) & (!g6) & (!g24) & (g3) & (g111)) + ((g42) & (!g45) & (g6) & (!g24) & (!g3) & (g111)) + ((g42) & (!g45) & (g6) & (!g24) & (g3) & (!g111)) + ((g42) & (!g45) & (g6) & (!g24) & (g3) & (g111)) + ((g42) & (!g45) & (g6) & (g24) & (g3) & (!g111)) + ((g42) & (!g45) & (g6) & (g24) & (g3) & (g111)) + ((g42) & (g45) & (g6) & (!g24) & (g3) & (!g111)) + ((g42) & (g45) & (g6) & (!g24) & (g3) & (g111)) + ((g42) & (g45) & (g6) & (g24) & (g3) & (!g111)) + ((g42) & (g45) & (g6) & (g24) & (g3) & (g111)));
	assign g124 = (((!g21) & (g2) & (g110)));
	assign g125 = (((!g12) & (!g123) & (!g105) & (!g86) & (!g124)) + ((!g12) & (!g123) & (!g105) & (g86) & (!g124)) + ((!g12) & (!g123) & (g105) & (!g86) & (!g124)) + ((!g12) & (!g123) & (g105) & (g86) & (!g124)) + ((!g12) & (g123) & (!g105) & (!g86) & (!g124)) + ((!g12) & (g123) & (g105) & (!g86) & (!g124)) + ((g12) & (!g123) & (g105) & (!g86) & (!g124)) + ((g12) & (!g123) & (g105) & (g86) & (!g124)) + ((g12) & (g123) & (g105) & (!g86) & (!g124)));
	assign g126 = (((!i_3_) & (!i_4_) & (!i_5_) & (!i_0_) & (!i_1_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (!i_0_) & (i_1_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (i_0_) & (i_1_)) + ((!i_3_) & (!i_4_) & (i_5_) & (!i_0_) & (!i_1_)) + ((!i_3_) & (!i_4_) & (i_5_) & (!i_0_) & (i_1_)) + ((!i_3_) & (!i_4_) & (i_5_) & (i_0_) & (i_1_)) + ((!i_3_) & (i_4_) & (!i_5_) & (!i_0_) & (!i_1_)) + ((!i_3_) & (i_4_) & (!i_5_) & (!i_0_) & (i_1_)) + ((!i_3_) & (i_4_) & (!i_5_) & (i_0_) & (!i_1_)) + ((!i_3_) & (i_4_) & (!i_5_) & (i_0_) & (i_1_)) + ((!i_3_) & (i_4_) & (i_5_) & (!i_0_) & (!i_1_)) + ((!i_3_) & (i_4_) & (i_5_) & (!i_0_) & (i_1_)) + ((!i_3_) & (i_4_) & (i_5_) & (i_0_) & (!i_1_)) + ((!i_3_) & (i_4_) & (i_5_) & (i_0_) & (i_1_)) + ((i_3_) & (!i_4_) & (!i_5_) & (!i_0_) & (!i_1_)) + ((i_3_) & (!i_4_) & (!i_5_) & (!i_0_) & (i_1_)) + ((i_3_) & (!i_4_) & (!i_5_) & (i_0_) & (!i_1_)) + ((i_3_) & (!i_4_) & (!i_5_) & (i_0_) & (i_1_)) + ((i_3_) & (!i_4_) & (i_5_) & (!i_0_) & (!i_1_)) + ((i_3_) & (!i_4_) & (i_5_) & (!i_0_) & (i_1_)) + ((i_3_) & (!i_4_) & (i_5_) & (i_0_) & (!i_1_)) + ((i_3_) & (!i_4_) & (i_5_) & (i_0_) & (i_1_)) + ((i_3_) & (i_4_) & (!i_5_) & (!i_0_) & (!i_1_)) + ((i_3_) & (i_4_) & (!i_5_) & (i_0_) & (!i_1_)) + ((i_3_) & (i_4_) & (!i_5_) & (i_0_) & (i_1_)) + ((i_3_) & (i_4_) & (i_5_) & (!i_0_) & (!i_1_)) + ((i_3_) & (i_4_) & (i_5_) & (!i_0_) & (i_1_)) + ((i_3_) & (i_4_) & (i_5_) & (i_0_) & (!i_1_)) + ((i_3_) & (i_4_) & (i_5_) & (i_0_) & (i_1_)));
	assign g140 = (((!g27) & (!g6) & (!g36) & (!g138) & (!g139)) + ((!g27) & (!g6) & (g36) & (!g138) & (!g139)) + ((!g27) & (g6) & (g36) & (!g138) & (!g139)) + ((g27) & (!g6) & (!g36) & (!g138) & (!g139)) + ((g27) & (!g6) & (g36) & (!g138) & (!g139)) + ((g27) & (g6) & (!g36) & (!g138) & (!g139)) + ((g27) & (g6) & (g36) & (!g138) & (!g139)));
	assign g145 = (((!i_6_) & (g137) & (!g51) & (g33) & (!g85)) + ((!i_6_) & (g137) & (!g51) & (g33) & (g85)) + ((!i_6_) & (g137) & (g51) & (!g33) & (g85)) + ((!i_6_) & (g137) & (g51) & (g33) & (!g85)) + ((!i_6_) & (g137) & (g51) & (g33) & (g85)) + ((i_6_) & (g137) & (g51) & (!g33) & (g85)) + ((i_6_) & (g137) & (g51) & (g33) & (g85)));
	assign g147 = (((!g37) & (!g38) & (!g110) & (!g145) & (!g146)) + ((!g37) & (!g38) & (g110) & (!g145) & (!g146)) + ((!g37) & (g38) & (!g110) & (!g145) & (!g146)) + ((!g37) & (g38) & (g110) & (!g145) & (!g146)) + ((g37) & (!g38) & (!g110) & (!g145) & (!g146)) + ((g37) & (g38) & (!g110) & (!g145) & (!g146)) + ((g37) & (g38) & (g110) & (!g145) & (!g146)));
	assign g149 = (((!g21) & (!g23) & (!g7) & (g100)) + ((!g21) & (!g23) & (g7) & (!g100)) + ((!g21) & (!g23) & (g7) & (g100)) + ((!g21) & (g23) & (g7) & (!g100)) + ((!g21) & (g23) & (g7) & (g100)) + ((g21) & (!g23) & (!g7) & (g100)) + ((g21) & (!g23) & (g7) & (g100)));
	assign g152 = (((!g6) & (!g77) & (!g148) & (!g149) & (g151)) + ((!g6) & (g77) & (!g148) & (!g149) & (g151)) + ((g6) & (!g77) & (!g148) & (!g149) & (g151)));
	assign g154 = (((g115) & (g119) & (g133) & (g144) & (g153)));
	assign g157 = (((!g47) & (!g75) & (!g155) & (!g156)) + ((!g47) & (g75) & (!g155) & (!g156)) + ((g47) & (!g75) & (!g155) & (!g156)));
	assign g160 = (((!g42) & (g12) & (g84) & (!g159)) + ((!g42) & (g12) & (g84) & (g159)) + ((g42) & (!g12) & (!g84) & (g159)) + ((g42) & (!g12) & (g84) & (g159)) + ((g42) & (g12) & (!g84) & (g159)) + ((g42) & (g12) & (g84) & (!g159)) + ((g42) & (g12) & (g84) & (g159)));
	assign g164 = (((!g2) & (!g158) & (!g160) & (!g162) & (!g163)) + ((!g2) & (g158) & (!g160) & (!g162) & (!g163)) + ((g2) & (!g158) & (!g160) & (!g162) & (!g163)));
	assign g165 = (((!g27) & (!g59) & (g60)));
	assign g166 = (((!i_5_) & (!g42) & (!g2) & (!g165)) + ((!i_5_) & (!g42) & (g2) & (!g165)) + ((!i_5_) & (g42) & (!g2) & (!g165)) + ((i_5_) & (!g42) & (!g2) & (!g165)) + ((i_5_) & (!g42) & (g2) & (!g165)) + ((i_5_) & (g42) & (!g2) & (!g165)) + ((i_5_) & (g42) & (g2) & (!g165)));
	assign g168 = (((!i_0_) & (!i_2_) & (g35) & (g75) & (!g167)) + ((!i_0_) & (!i_2_) & (g35) & (g75) & (g167)) + ((!i_0_) & (i_2_) & (g35) & (g75) & (!g167)) + ((!i_0_) & (i_2_) & (g35) & (g75) & (g167)) + ((i_0_) & (!i_2_) & (g35) & (g75) & (!g167)) + ((i_0_) & (!i_2_) & (g35) & (g75) & (g167)) + ((i_0_) & (i_2_) & (!g35) & (!g75) & (g167)) + ((i_0_) & (i_2_) & (!g35) & (g75) & (g167)) + ((i_0_) & (i_2_) & (g35) & (!g75) & (g167)) + ((i_0_) & (i_2_) & (g35) & (g75) & (!g167)) + ((i_0_) & (i_2_) & (g35) & (g75) & (g167)));
	assign g170 = (((i_3_) & (!i_5_) & (!g25) & (g12)));
	assign g173 = (((g127) & (!i_2_) & (g8) & (!g45) & (!g12)) + ((g127) & (!i_2_) & (g8) & (!g45) & (g12)) + ((g127) & (i_2_) & (!g8) & (!g45) & (g12)) + ((g127) & (i_2_) & (g8) & (!g45) & (g12)));
	assign g174 = (((!g11) & (!g8) & (g29) & (!g91)) + ((!g11) & (!g8) & (g29) & (g91)) + ((!g11) & (g8) & (!g29) & (g91)) + ((!g11) & (g8) & (g29) & (!g91)) + ((!g11) & (g8) & (g29) & (g91)) + ((g11) & (g8) & (!g29) & (g91)) + ((g11) & (g8) & (g29) & (g91)));
	assign g175 = (((!g25) & (!g45) & (!g22) & (g6)) + ((!g25) & (!g45) & (g22) & (!g6)) + ((!g25) & (!g45) & (g22) & (g6)) + ((!g25) & (g45) & (g22) & (!g6)) + ((!g25) & (g45) & (g22) & (g6)));
	assign g178 = (((!g11) & (!g9) & (!g169) & (g172) & (g177)) + ((g11) & (!g9) & (!g169) & (g172) & (g177)) + ((g11) & (g9) & (!g169) & (g172) & (g177)));
	assign g179 = (((!g35) & (!g21) & (g12) & (!g24) & (!g26)) + ((!g35) & (!g21) & (g12) & (!g24) & (g26)) + ((g35) & (!g21) & (!g12) & (!g24) & (g26)) + ((g35) & (!g21) & (!g12) & (g24) & (g26)) + ((g35) & (!g21) & (g12) & (!g24) & (!g26)) + ((g35) & (!g21) & (g12) & (!g24) & (g26)) + ((g35) & (!g21) & (g12) & (g24) & (g26)) + ((g35) & (g21) & (!g12) & (!g24) & (g26)) + ((g35) & (g21) & (!g12) & (g24) & (g26)) + ((g35) & (g21) & (g12) & (!g24) & (g26)) + ((g35) & (g21) & (g12) & (g24) & (g26)));
	assign g186 = (((!g45) & (!g48) & (g2) & (!g24) & (g184)) + ((!g45) & (!g48) & (g2) & (g24) & (g184)) + ((!g45) & (g48) & (!g2) & (!g24) & (!g184)) + ((!g45) & (g48) & (!g2) & (!g24) & (g184)) + ((!g45) & (g48) & (g2) & (!g24) & (!g184)) + ((!g45) & (g48) & (g2) & (!g24) & (g184)) + ((!g45) & (g48) & (g2) & (g24) & (g184)) + ((g45) & (!g48) & (g2) & (!g24) & (g184)) + ((g45) & (!g48) & (g2) & (g24) & (g184)) + ((g45) & (g48) & (g2) & (!g24) & (g184)) + ((g45) & (g48) & (g2) & (g24) & (g184)));
	assign g187 = (((!i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (i_6_) & (i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (!i_5_) & (i_6_) & (i_7_) & (i_8_)) + ((!i_3_) & (!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (!i_4_) & (i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (i_5_) & (!i_6_) & (i_7_) & (i_8_)) + ((!i_3_) & (!i_4_) & (i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (i_5_) & (i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (!i_4_) & (i_5_) & (i_6_) & (i_7_) & (!i_8_)) + ((!i_3_) & (!i_4_) & (i_5_) & (i_6_) & (i_7_) & (i_8_)) + ((!i_3_) & (i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_8_)) + ((!i_3_) & (i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((!i_3_) & (i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (i_8_)) + ((!i_3_) & (i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((!i_3_) & (i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (i_4_) & (!i_5_) & (i_6_) & (i_7_) & (!i_8_)) + ((!i_3_) & (i_4_) & (!i_5_) & (i_6_) & (i_7_) & (i_8_)) + ((!i_3_) & (i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (i_4_) & (i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((!i_3_) & (i_4_) & (i_5_) & (!i_6_) & (i_7_) & (i_8_)) + ((!i_3_) & (i_4_) & (i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((!i_3_) & (i_4_) & (i_5_) & (i_6_) & (!i_7_) & (i_8_)) + ((!i_3_) & (i_4_) & (i_5_) & (i_6_) & (i_7_) & (!i_8_)) + ((!i_3_) & (i_4_) & (i_5_) & (i_6_) & (i_7_) & (i_8_)) + ((i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_8_)) + ((i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (i_8_)) + ((i_3_) & (!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((i_3_) & (!i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (i_8_)) + ((i_3_) & (!i_4_) & (!i_5_) & (i_6_) & (i_7_) & (!i_8_)) + ((i_3_) & (!i_4_) & (!i_5_) & (i_6_) & (i_7_) & (i_8_)) + ((i_3_) & (!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((i_3_) & (!i_4_) & (i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((i_3_) & (!i_4_) & (i_5_) & (!i_6_) & (i_7_) & (i_8_)) + ((i_3_) & (!i_4_) & (i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((i_3_) & (!i_4_) & (i_5_) & (i_6_) & (!i_7_) & (i_8_)) + ((i_3_) & (!i_4_) & (i_5_) & (i_6_) & (i_7_) & (!i_8_)) + ((i_3_) & (!i_4_) & (i_5_) & (i_6_) & (i_7_) & (i_8_)) + ((i_3_) & (i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (!i_8_)) + ((i_3_) & (i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((i_3_) & (i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((i_3_) & (i_4_) & (!i_5_) & (i_6_) & (!i_7_) & (i_8_)) + ((i_3_) & (i_4_) & (!i_5_) & (i_6_) & (i_7_) & (!i_8_)) + ((i_3_) & (i_4_) & (!i_5_) & (i_6_) & (i_7_) & (i_8_)) + ((i_3_) & (i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((i_3_) & (i_4_) & (i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((i_3_) & (i_4_) & (i_5_) & (!i_6_) & (i_7_) & (i_8_)) + ((i_3_) & (i_4_) & (i_5_) & (i_6_) & (!i_7_) & (!i_8_)) + ((i_3_) & (i_4_) & (i_5_) & (i_6_) & (!i_7_) & (i_8_)) + ((i_3_) & (i_4_) & (i_5_) & (i_6_) & (i_7_) & (!i_8_)) + ((i_3_) & (i_4_) & (i_5_) & (i_6_) & (i_7_) & (i_8_)));
	assign g188 = (((i_3_) & (!i_5_) & (g35) & (g42)));
	assign g193 = (((!g23) & (!g3) & (!g7) & (g181)) + ((!g23) & (!g3) & (g7) & (g181)) + ((!g23) & (g3) & (!g7) & (g181)) + ((!g23) & (g3) & (g7) & (!g181)) + ((!g23) & (g3) & (g7) & (g181)) + ((g23) & (g3) & (g7) & (!g181)) + ((g23) & (g3) & (g7) & (g181)));
	assign g195 = (((!g8) & (!g13) & (!g181) & (g194)) + ((!g8) & (!g13) & (g181) & (g194)) + ((g8) & (!g13) & (!g181) & (g194)) + ((g8) & (!g13) & (g181) & (!g194)) + ((g8) & (!g13) & (g181) & (g194)) + ((g8) & (g13) & (g181) & (!g194)) + ((g8) & (g13) & (g181) & (g194)));
	assign g200 = (((!g27) & (!g45) & (!g23) & (!g36) & (!g121)) + ((!g27) & (!g45) & (!g23) & (!g36) & (g121)) + ((!g27) & (!g45) & (!g23) & (g36) & (!g121)) + ((!g27) & (!g45) & (!g23) & (g36) & (g121)) + ((!g27) & (!g45) & (g23) & (!g36) & (g121)) + ((!g27) & (g45) & (!g23) & (!g36) & (g121)) + ((!g27) & (g45) & (g23) & (!g36) & (g121)) + ((g27) & (!g45) & (!g23) & (!g36) & (g121)) + ((g27) & (!g45) & (g23) & (!g36) & (g121)) + ((g27) & (g45) & (!g23) & (!g36) & (g121)) + ((g27) & (g45) & (g23) & (!g36) & (g121)));
	assign g202 = (((!g45) & (!g37) & (!g13) & (!g201)) + ((!g45) & (!g37) & (g13) & (!g201)) + ((!g45) & (g37) & (g13) & (!g201)) + ((g45) & (!g37) & (!g13) & (!g201)) + ((g45) & (!g37) & (g13) & (!g201)) + ((g45) & (g37) & (!g13) & (!g201)) + ((g45) & (g37) & (g13) & (!g201)));
	assign g204 = (((!i_6_) & (!i_8_) & (g32) & (!g105) & (g141)) + ((!i_6_) & (!i_8_) & (g32) & (g105) & (g141)) + ((!i_6_) & (i_8_) & (g32) & (!g105) & (g141)) + ((!i_6_) & (i_8_) & (g32) & (g105) & (g141)) + ((i_6_) & (!i_8_) & (g32) & (!g105) & (g141)) + ((i_6_) & (!i_8_) & (g32) & (g105) & (g141)) + ((i_6_) & (i_8_) & (!g32) & (!g105) & (!g141)) + ((i_6_) & (i_8_) & (!g32) & (!g105) & (g141)) + ((i_6_) & (i_8_) & (g32) & (!g105) & (!g141)) + ((i_6_) & (i_8_) & (g32) & (!g105) & (g141)) + ((i_6_) & (i_8_) & (g32) & (g105) & (g141)));
	assign g206 = (((!g150) & (!g200) & (g202) & (!g203) & (g205)));
	assign g208 = (((!i_6_) & (!g42) & (g46) & (g47) & (!g38)) + ((!i_6_) & (!g42) & (g46) & (g47) & (g38)) + ((!i_6_) & (g42) & (g46) & (g47) & (!g38)) + ((!i_6_) & (g42) & (g46) & (g47) & (g38)) + ((i_6_) & (g42) & (!g46) & (g47) & (!g38)) + ((i_6_) & (g42) & (g46) & (g47) & (!g38)));
	assign g211 = (((!g1) & (!g47) & (!g64) & (!g207) & (g210)) + ((!g1) & (!g47) & (g64) & (!g207) & (g210)) + ((!g1) & (g47) & (!g64) & (!g207) & (g210)) + ((g1) & (!g47) & (!g64) & (!g207) & (g210)) + ((g1) & (!g47) & (g64) & (!g207) & (g210)) + ((g1) & (g47) & (!g64) & (!g207) & (g210)) + ((g1) & (g47) & (g64) & (!g207) & (g210)));
	assign g215 = (((!i_4_) & (!i_5_) & (!g6) & (!g13) & (g214)) + ((!i_4_) & (!i_5_) & (!g6) & (g13) & (g214)) + ((!i_4_) & (!i_5_) & (g6) & (!g13) & (g214)) + ((!i_4_) & (!i_5_) & (g6) & (g13) & (g214)) + ((!i_4_) & (i_5_) & (!g6) & (!g13) & (g214)) + ((!i_4_) & (i_5_) & (!g6) & (g13) & (g214)) + ((!i_4_) & (i_5_) & (g6) & (!g13) & (g214)) + ((!i_4_) & (i_5_) & (g6) & (g13) & (g214)) + ((i_4_) & (!i_5_) & (!g6) & (!g13) & (g214)) + ((i_4_) & (!i_5_) & (!g6) & (g13) & (g214)) + ((i_4_) & (!i_5_) & (g6) & (!g13) & (g214)) + ((i_4_) & (!i_5_) & (g6) & (g13) & (g214)) + ((i_4_) & (i_5_) & (!g6) & (!g13) & (g214)) + ((i_4_) & (i_5_) & (!g6) & (g13) & (g214)) + ((i_4_) & (i_5_) & (g6) & (g13) & (g214)));
	assign g216 = (((!i_1_) & (!g135) & (!g212) & (g215)) + ((i_1_) & (!g135) & (!g212) & (g215)) + ((i_1_) & (g135) & (!g212) & (g215)));
	assign g218 = (((g42) & (g217)));
	assign g224 = (((!i_7_) & (!g218) & (!g220) & (g222) & (g223)) + ((i_7_) & (!g218) & (!g220) & (g222) & (g223)) + ((i_7_) & (g218) & (!g220) & (g222) & (g223)));
	assign g226 = (((!g63) & (g41) & (!g1) & (!g36) & (!g225)) + ((!g63) & (g41) & (!g1) & (!g36) & (g225)) + ((!g63) & (g41) & (g1) & (!g36) & (!g225)) + ((!g63) & (g41) & (g1) & (!g36) & (g225)) + ((g63) & (!g41) & (!g1) & (!g36) & (g225)) + ((g63) & (!g41) & (!g1) & (g36) & (g225)) + ((g63) & (g41) & (!g1) & (!g36) & (!g225)) + ((g63) & (g41) & (!g1) & (!g36) & (g225)) + ((g63) & (g41) & (!g1) & (g36) & (g225)) + ((g63) & (g41) & (g1) & (!g36) & (!g225)) + ((g63) & (g41) & (g1) & (!g36) & (g225)));
	assign g228 = (((!g186) & (!g226) & (!g227)));
	assign g229 = (((!g23) & (!g71) & (g161)) + ((!g23) & (g71) & (!g161)) + ((!g23) & (g71) & (g161)));
	assign g234 = (((!g30) & (g216) & (g224) & (g228) & (g233)));
	assign g236 = (((!g6) & (!g73) & (!g49) & (!g60) & (!g235)) + ((!g6) & (!g73) & (!g49) & (g60) & (!g235)) + ((!g6) & (!g73) & (g49) & (!g60) & (!g235)) + ((!g6) & (g73) & (!g49) & (!g60) & (!g235)) + ((!g6) & (g73) & (!g49) & (g60) & (!g235)) + ((!g6) & (g73) & (g49) & (!g60) & (!g235)) + ((g6) & (!g73) & (!g49) & (!g60) & (!g235)) + ((g6) & (!g73) & (!g49) & (g60) & (!g235)) + ((g6) & (!g73) & (g49) & (!g60) & (!g235)));
	assign g239 = (((!g11) & (!g45) & (!g2) & (!g23) & (!g13)) + ((!g11) & (!g45) & (g2) & (!g23) & (!g13)) + ((!g11) & (!g45) & (g2) & (g23) & (!g13)) + ((!g11) & (g45) & (!g2) & (!g23) & (!g13)) + ((!g11) & (g45) & (g2) & (!g23) & (!g13)) + ((g11) & (!g45) & (g2) & (!g23) & (!g13)) + ((g11) & (!g45) & (g2) & (g23) & (!g13)));
	assign g242 = (((!g6) & (!g88) & (!g238) & (g241)) + ((!g6) & (g88) & (!g238) & (g241)) + ((g6) & (!g88) & (!g238) & (g241)));
	assign g244 = (((g63) & (g51) & (g134)));
	assign g246 = (((!i_6_) & (!i_8_) & (!g243) & (g245)) + ((!i_6_) & (!i_8_) & (g243) & (g245)) + ((!i_6_) & (i_8_) & (!g243) & (g245)) + ((i_6_) & (!i_8_) & (!g243) & (g245)) + ((i_6_) & (!i_8_) & (g243) & (g245)) + ((i_6_) & (i_8_) & (!g243) & (g245)) + ((i_6_) & (i_8_) & (g243) & (g245)));
	assign g247 = (((!g35) & (!g42) & (!g25) & (!g23) & (g3)) + ((!g35) & (g42) & (!g25) & (!g23) & (g3)) + ((g35) & (!g42) & (!g25) & (!g23) & (g3)) + ((g35) & (g42) & (!g25) & (!g23) & (g3)) + ((g35) & (g42) & (!g25) & (g23) & (g3)) + ((g35) & (g42) & (g25) & (!g23) & (g3)) + ((g35) & (g42) & (g25) & (g23) & (g3)));
	assign g249 = (((!g21) & (!g8) & (!g25) & (!g247) & (!g248)) + ((!g21) & (!g8) & (g25) & (!g247) & (!g248)) + ((!g21) & (g8) & (g25) & (!g247) & (!g248)) + ((g21) & (!g8) & (!g25) & (!g247) & (!g248)) + ((g21) & (!g8) & (g25) & (!g247) & (!g248)) + ((g21) & (g8) & (!g25) & (!g247) & (!g248)) + ((g21) & (g8) & (g25) & (!g247) & (!g248)));
	assign g251 = (((!i_3_) & (!i_0_) & (!i_1_) & (!g219) & (!g250)) + ((!i_3_) & (!i_0_) & (!i_1_) & (g219) & (!g250)) + ((!i_3_) & (!i_0_) & (i_1_) & (!g219) & (!g250)) + ((!i_3_) & (i_0_) & (!i_1_) & (!g219) & (!g250)) + ((!i_3_) & (i_0_) & (!i_1_) & (g219) & (!g250)) + ((!i_3_) & (i_0_) & (i_1_) & (!g219) & (!g250)) + ((!i_3_) & (i_0_) & (i_1_) & (g219) & (!g250)) + ((i_3_) & (!i_0_) & (!i_1_) & (!g219) & (!g250)) + ((i_3_) & (!i_0_) & (!i_1_) & (g219) & (!g250)) + ((i_3_) & (!i_0_) & (i_1_) & (!g219) & (!g250)) + ((i_3_) & (!i_0_) & (i_1_) & (g219) & (!g250)) + ((i_3_) & (i_0_) & (!i_1_) & (!g219) & (!g250)) + ((i_3_) & (i_0_) & (!i_1_) & (g219) & (!g250)) + ((i_3_) & (i_0_) & (i_1_) & (!g219) & (!g250)) + ((i_3_) & (i_0_) & (i_1_) & (g219) & (!g250)));
	assign g254 = (((!g127) & (!g6) & (!g5) & (g251) & (g253)) + ((!g127) & (!g6) & (g5) & (g251) & (g253)) + ((!g127) & (g6) & (!g5) & (g251) & (g253)) + ((!g127) & (g6) & (g5) & (g251) & (g253)) + ((g127) & (!g6) & (!g5) & (g251) & (g253)) + ((g127) & (!g6) & (g5) & (g251) & (g253)) + ((g127) & (g6) & (!g5) & (g251) & (g253)));
	assign g255 = (((!g14) & (!g1) & (g12) & (g3) & (!g225)) + ((!g14) & (!g1) & (g12) & (g3) & (g225)) + ((g14) & (!g1) & (!g12) & (!g3) & (g225)) + ((g14) & (!g1) & (!g12) & (g3) & (g225)) + ((g14) & (!g1) & (g12) & (!g3) & (g225)) + ((g14) & (!g1) & (g12) & (g3) & (!g225)) + ((g14) & (!g1) & (g12) & (g3) & (g225)));
	assign g256 = (((!g25) & (g120) & (!g23)));
	assign g257 = (((!g8) & (!g1) & (!g22) & (!g105) & (!g256)) + ((!g8) & (!g1) & (!g22) & (g105) & (!g256)) + ((!g8) & (g1) & (!g22) & (!g105) & (!g256)) + ((!g8) & (g1) & (!g22) & (g105) & (!g256)) + ((!g8) & (g1) & (g22) & (!g105) & (!g256)) + ((!g8) & (g1) & (g22) & (g105) & (!g256)) + ((g8) & (!g1) & (!g22) & (g105) & (!g256)) + ((g8) & (g1) & (!g22) & (g105) & (!g256)) + ((g8) & (g1) & (g22) & (g105) & (!g256)));
	assign g264 = (((!g11) & (!g42) & (!g23) & (!g13) & (!g60) & (!g38)) + ((!g11) & (!g42) & (!g23) & (!g13) & (g60) & (!g38)) + ((!g11) & (g42) & (!g23) & (!g13) & (!g60) & (!g38)) + ((!g11) & (g42) & (!g23) & (!g13) & (g60) & (!g38)) + ((!g11) & (g42) & (!g23) & (!g13) & (g60) & (g38)) + ((!g11) & (g42) & (!g23) & (g13) & (g60) & (!g38)) + ((!g11) & (g42) & (!g23) & (g13) & (g60) & (g38)) + ((!g11) & (g42) & (g23) & (!g13) & (g60) & (!g38)) + ((!g11) & (g42) & (g23) & (!g13) & (g60) & (g38)) + ((!g11) & (g42) & (g23) & (g13) & (g60) & (!g38)) + ((!g11) & (g42) & (g23) & (g13) & (g60) & (g38)) + ((g11) & (!g42) & (!g23) & (!g13) & (!g60) & (!g38)) + ((g11) & (!g42) & (!g23) & (!g13) & (g60) & (!g38)) + ((g11) & (g42) & (!g23) & (!g13) & (!g60) & (!g38)) + ((g11) & (g42) & (!g23) & (!g13) & (g60) & (!g38)));
	assign g266 = (((!g11) & (!g12) & (!g71) & (g265)) + ((!g11) & (!g12) & (g71) & (g265)) + ((!g11) & (g12) & (!g71) & (g265)) + ((!g11) & (g12) & (g71) & (!g265)) + ((!g11) & (g12) & (g71) & (g265)) + ((g11) & (g12) & (g71) & (!g265)) + ((g11) & (g12) & (g71) & (g265)));
	assign g267 = (((!g27) & (!g35) & (!g36) & (!g110) & (g194)) + ((!g27) & (!g35) & (!g36) & (g110) & (g194)) + ((!g27) & (!g35) & (g36) & (!g110) & (g194)) + ((!g27) & (!g35) & (g36) & (g110) & (g194)) + ((!g27) & (g35) & (!g36) & (!g110) & (g194)) + ((!g27) & (g35) & (!g36) & (g110) & (!g194)) + ((!g27) & (g35) & (!g36) & (g110) & (g194)) + ((!g27) & (g35) & (g36) & (!g110) & (g194)) + ((!g27) & (g35) & (g36) & (g110) & (g194)) + ((g27) & (g35) & (!g36) & (g110) & (!g194)) + ((g27) & (g35) & (!g36) & (g110) & (g194)));
	assign g268 = (((!g24) & (g225)));
	assign g274 = (((!g264) & (!g266) & (!g267) & (g215) & (g273)));
	assign g275 = (((!g27) & (i_7_) & (!i_8_) & (!g36) & (!g100)) + ((!g27) & (i_7_) & (!i_8_) & (!g36) & (g100)) + ((!g27) & (i_7_) & (i_8_) & (!g36) & (g100)) + ((!g27) & (i_7_) & (i_8_) & (g36) & (g100)) + ((g27) & (i_7_) & (i_8_) & (!g36) & (g100)) + ((g27) & (i_7_) & (i_8_) & (g36) & (g100)));
	assign g276 = (((!g28) & (!g42) & (!g23) & (!g3) & (g91)) + ((!g28) & (!g42) & (!g23) & (g3) & (g91)) + ((!g28) & (g42) & (!g23) & (!g3) & (g91)) + ((!g28) & (g42) & (!g23) & (g3) & (g91)) + ((g28) & (!g42) & (!g23) & (!g3) & (g91)) + ((g28) & (!g42) & (!g23) & (g3) & (g91)) + ((g28) & (g42) & (!g23) & (!g3) & (g91)) + ((g28) & (g42) & (!g23) & (g3) & (!g91)) + ((g28) & (g42) & (!g23) & (g3) & (g91)) + ((g28) & (g42) & (g23) & (g3) & (!g91)) + ((g28) & (g42) & (g23) & (g3) & (g91)));
	assign g277 = (((!g11) & (!g8) & (g12) & (!g13) & (!g184)) + ((!g11) & (!g8) & (g12) & (!g13) & (g184)) + ((!g11) & (g8) & (!g12) & (!g13) & (g184)) + ((!g11) & (g8) & (!g12) & (g13) & (g184)) + ((!g11) & (g8) & (g12) & (!g13) & (!g184)) + ((!g11) & (g8) & (g12) & (!g13) & (g184)) + ((!g11) & (g8) & (g12) & (g13) & (g184)) + ((g11) & (g8) & (!g12) & (!g13) & (g184)) + ((g11) & (g8) & (!g12) & (g13) & (g184)) + ((g11) & (g8) & (g12) & (!g13) & (g184)) + ((g11) & (g8) & (g12) & (g13) & (g184)));
	assign g278 = (((g35) & (!g46) & (g158)) + ((g35) & (g46) & (!g158)) + ((g35) & (g46) & (g158)));
	assign g279 = (((!g38) & (!g94) & (g265) & (!g167)) + ((!g38) & (!g94) & (g265) & (g167)) + ((!g38) & (g94) & (!g265) & (g167)) + ((!g38) & (g94) & (g265) & (!g167)) + ((!g38) & (g94) & (g265) & (g167)) + ((g38) & (g94) & (!g265) & (g167)) + ((g38) & (g94) & (g265) & (g167)));
	assign g283 = (((!i_0_) & (!g135) & (!g275) & (!g276) & (g282)) + ((!i_0_) & (g135) & (!g275) & (!g276) & (g282)) + ((i_0_) & (!g135) & (!g275) & (!g276) & (g282)));
	assign g285 = (((!i_6_) & (!i_8_) & (!g1) & (g32)));
	assign g287 = (((!g25) & (!g194) & (!g212) & (!g285) & (g286)) + ((g25) & (!g194) & (!g212) & (!g285) & (g286)) + ((g25) & (g194) & (!g212) & (!g285) & (g286)));
	assign g289 = (((!g13) & (!g123) & (!g284) & (g287) & (!g288)) + ((g13) & (!g123) & (!g284) & (g287) & (!g288)) + ((g13) & (g123) & (!g284) & (g287) & (!g288)));
	assign g291 = (((!g48) & (!g181) & (!g244) & (!g290)) + ((!g48) & (g181) & (!g244) & (!g290)) + ((g48) & (!g181) & (!g244) & (!g290)));
	assign g292 = (((!g27) & (i_6_) & (!i_8_) & (!g21)));
	assign g293 = (((!g27) & (!g35) & (!g45) & (g6) & (!g84)) + ((!g27) & (!g35) & (!g45) & (g6) & (g84)) + ((!g27) & (g35) & (!g45) & (!g6) & (g84)) + ((!g27) & (g35) & (!g45) & (g6) & (!g84)) + ((!g27) & (g35) & (!g45) & (g6) & (g84)) + ((!g27) & (g35) & (g45) & (!g6) & (g84)) + ((!g27) & (g35) & (g45) & (g6) & (g84)) + ((g27) & (g35) & (!g45) & (!g6) & (g84)) + ((g27) & (g35) & (!g45) & (g6) & (g84)) + ((g27) & (g35) & (g45) & (!g6) & (g84)) + ((g27) & (g35) & (g45) & (g6) & (g84)));
	assign g300 = (((g164) & (g283) & (g289) & (g291) & (g299)));
	assign g301 = (((!i_6_) & (g137) & (!g77) & (!g13) & (g64)) + ((!i_6_) & (g137) & (g77) & (!g13) & (!g64)) + ((!i_6_) & (g137) & (g77) & (!g13) & (g64)) + ((!i_6_) & (g137) & (g77) & (g13) & (!g64)) + ((!i_6_) & (g137) & (g77) & (g13) & (g64)) + ((i_6_) & (g137) & (!g77) & (!g13) & (g64)) + ((i_6_) & (g137) & (g77) & (!g13) & (g64)));
	assign g307 = (((!g11) & (!g67) & (!g302) & (g303) & (g306)) + ((g11) & (!g67) & (!g302) & (g303) & (g306)) + ((g11) & (g67) & (!g302) & (g303) & (g306)));
	assign g310 = (((!i_6_) & (!i_7_) & (!g129) & (!g309)) + ((!i_6_) & (!i_7_) & (g129) & (!g309)) + ((!i_6_) & (i_7_) & (!g129) & (!g309)) + ((!i_6_) & (i_7_) & (g129) & (!g309)) + ((i_6_) & (!i_7_) & (!g129) & (!g309)) + ((i_6_) & (i_7_) & (!g129) & (!g309)) + ((i_6_) & (i_7_) & (g129) & (!g309)));
	assign g312 = (((!i_3_) & (!i_4_) & (!g28) & (!g24) & (!g311)) + ((!i_3_) & (!i_4_) & (!g28) & (g24) & (!g311)) + ((!i_3_) & (!i_4_) & (g28) & (!g24) & (!g311)) + ((!i_3_) & (!i_4_) & (g28) & (g24) & (!g311)) + ((!i_3_) & (i_4_) & (!g28) & (!g24) & (!g311)) + ((!i_3_) & (i_4_) & (!g28) & (g24) & (!g311)) + ((!i_3_) & (i_4_) & (g28) & (!g24) & (!g311)) + ((!i_3_) & (i_4_) & (g28) & (g24) & (!g311)) + ((i_3_) & (!i_4_) & (!g28) & (!g24) & (!g311)) + ((i_3_) & (!i_4_) & (!g28) & (g24) & (!g311)) + ((i_3_) & (!i_4_) & (g28) & (g24) & (!g311)) + ((i_3_) & (i_4_) & (!g28) & (!g24) & (!g311)) + ((i_3_) & (i_4_) & (!g28) & (g24) & (!g311)) + ((i_3_) & (i_4_) & (g28) & (!g24) & (!g311)) + ((i_3_) & (i_4_) & (g28) & (g24) & (!g311)));
	assign g313 = (((!g25) & (!g12) & (!g32) & (g9) & (g116)) + ((!g25) & (!g12) & (g32) & (g9) & (g116)) + ((!g25) & (g12) & (!g32) & (g9) & (g116)) + ((!g25) & (g12) & (g32) & (!g9) & (!g116)) + ((!g25) & (g12) & (g32) & (!g9) & (g116)) + ((!g25) & (g12) & (g32) & (g9) & (!g116)) + ((!g25) & (g12) & (g32) & (g9) & (g116)) + ((g25) & (!g12) & (!g32) & (g9) & (g116)) + ((g25) & (!g12) & (g32) & (g9) & (g116)) + ((g25) & (g12) & (!g32) & (g9) & (g116)) + ((g25) & (g12) & (g32) & (g9) & (g116)));
	assign g314 = (((!g11) & (!g48) & (!g24) & (!g32) & (g9)) + ((!g11) & (!g48) & (!g24) & (g32) & (g9)) + ((!g11) & (!g48) & (g24) & (!g32) & (g9)) + ((!g11) & (!g48) & (g24) & (g32) & (g9)) + ((!g11) & (g48) & (!g24) & (!g32) & (g9)) + ((!g11) & (g48) & (!g24) & (g32) & (!g9)) + ((!g11) & (g48) & (!g24) & (g32) & (g9)) + ((!g11) & (g48) & (g24) & (!g32) & (g9)) + ((!g11) & (g48) & (g24) & (g32) & (g9)) + ((g11) & (g48) & (!g24) & (g32) & (!g9)) + ((g11) & (g48) & (!g24) & (g32) & (g9)));
	assign g315 = (((!g1) & (g32) & (g37)));
	assign g323 = (((!g264) & (!g279) & (g596) & (!g321) & (!g322)));
	assign g327 = (((!g35) & (!g181) & (!g276) & (!g324) & (g326)) + ((!g35) & (g181) & (!g276) & (!g324) & (g326)) + ((g35) & (!g181) & (!g276) & (!g324) & (g326)));
	assign g330 = (((!g32) & (!g29) & (!g193) & (!g328) & (!g329)) + ((!g32) & (g29) & (!g193) & (!g328) & (!g329)) + ((g32) & (!g29) & (!g193) & (!g328) & (!g329)));
	assign g332 = (((!g45) & (!g2) & (!g49) & (!g7) & (!g331)) + ((!g45) & (!g2) & (g49) & (!g7) & (!g331)) + ((!g45) & (g2) & (!g49) & (!g7) & (!g331)) + ((g45) & (!g2) & (!g49) & (!g7) & (!g331)) + ((g45) & (!g2) & (!g49) & (g7) & (!g331)) + ((g45) & (!g2) & (g49) & (!g7) & (!g331)) + ((g45) & (!g2) & (g49) & (g7) & (!g331)) + ((g45) & (g2) & (!g49) & (!g7) & (!g331)) + ((g45) & (g2) & (!g49) & (g7) & (!g331)));
	assign g334 = (((i_3_) & (!g27) & (!i_6_) & (g333)));
	assign g341 = (((g119) & (g206) & (g327) & (g330) & (g340)));
	assign g343 = (((!g27) & (!g23) & (g36) & (!g285)) + ((!g27) & (g23) & (!g36) & (!g285)) + ((!g27) & (g23) & (g36) & (!g285)) + ((g27) & (!g23) & (!g36) & (!g285)) + ((g27) & (!g23) & (g36) & (!g285)) + ((g27) & (g23) & (!g36) & (!g285)) + ((g27) & (g23) & (g36) & (!g285)));
	assign g344 = (((!g21) & (!g6) & (!g23) & (!g24) & (!g129)) + ((!g21) & (!g6) & (!g23) & (!g24) & (g129)) + ((!g21) & (g6) & (!g23) & (!g24) & (!g129)) + ((!g21) & (g6) & (!g23) & (!g24) & (g129)) + ((!g21) & (g6) & (!g23) & (g24) & (g129)) + ((!g21) & (g6) & (g23) & (!g24) & (g129)) + ((!g21) & (g6) & (g23) & (g24) & (g129)) + ((g21) & (g6) & (!g23) & (!g24) & (g129)) + ((g21) & (g6) & (!g23) & (g24) & (g129)) + ((g21) & (g6) & (g23) & (!g24) & (g129)) + ((g21) & (g6) & (g23) & (g24) & (g129)));
	assign g346 = (((!g28) & (!g42) & (!g38) & (g110) & (g159) & (!g345)) + ((!g28) & (!g42) & (!g38) & (g110) & (g159) & (g345)) + ((!g28) & (!g42) & (g38) & (g110) & (g159) & (!g345)) + ((!g28) & (!g42) & (g38) & (g110) & (g159) & (g345)) + ((!g28) & (g42) & (!g38) & (!g110) & (!g159) & (g345)) + ((!g28) & (g42) & (!g38) & (!g110) & (g159) & (g345)) + ((!g28) & (g42) & (!g38) & (g110) & (!g159) & (g345)) + ((!g28) & (g42) & (!g38) & (g110) & (g159) & (!g345)) + ((!g28) & (g42) & (!g38) & (g110) & (g159) & (g345)) + ((!g28) & (g42) & (g38) & (!g110) & (!g159) & (g345)) + ((!g28) & (g42) & (g38) & (!g110) & (g159) & (g345)) + ((!g28) & (g42) & (g38) & (g110) & (!g159) & (g345)) + ((!g28) & (g42) & (g38) & (g110) & (g159) & (!g345)) + ((!g28) & (g42) & (g38) & (g110) & (g159) & (g345)) + ((g28) & (!g42) & (!g38) & (g110) & (!g159) & (!g345)) + ((g28) & (!g42) & (!g38) & (g110) & (!g159) & (g345)) + ((g28) & (!g42) & (!g38) & (g110) & (g159) & (!g345)) + ((g28) & (!g42) & (!g38) & (g110) & (g159) & (g345)) + ((g28) & (!g42) & (g38) & (g110) & (g159) & (!g345)) + ((g28) & (!g42) & (g38) & (g110) & (g159) & (g345)) + ((g28) & (g42) & (!g38) & (!g110) & (!g159) & (g345)) + ((g28) & (g42) & (!g38) & (!g110) & (g159) & (g345)) + ((g28) & (g42) & (!g38) & (g110) & (!g159) & (!g345)) + ((g28) & (g42) & (!g38) & (g110) & (!g159) & (g345)) + ((g28) & (g42) & (!g38) & (g110) & (g159) & (!g345)) + ((g28) & (g42) & (!g38) & (g110) & (g159) & (g345)) + ((g28) & (g42) & (g38) & (!g110) & (!g159) & (g345)) + ((g28) & (g42) & (g38) & (!g110) & (g159) & (g345)) + ((g28) & (g42) & (g38) & (g110) & (!g159) & (g345)) + ((g28) & (g42) & (g38) & (g110) & (g159) & (!g345)) + ((g28) & (g42) & (g38) & (g110) & (g159) & (g345)));
	assign g352 = (((!i_3_) & (!i_0_) & (i_1_) & (!g351)));
	assign g358 = (((!i_6_) & (!i_7_) & (!g75) & (!g357)) + ((!i_6_) & (!i_7_) & (g75) & (!g357)) + ((!i_6_) & (i_7_) & (!g75) & (!g357)) + ((!i_6_) & (i_7_) & (g75) & (!g357)) + ((i_6_) & (!i_7_) & (!g75) & (!g357)) + ((i_6_) & (i_7_) & (!g75) & (!g357)) + ((i_6_) & (i_7_) & (g75) & (!g357)));
	assign g363 = (((i_4_) & (i_5_) & (!g23) & (g110)));
	assign g364 = (((!g21) & (g6) & (!g24)));
	assign g367 = (((g202) & (g358) & (!g360) & (g362) & (g366)));
	assign g368 = (((!g11) & (!g41) & (g28) & (g70)) + ((!g11) & (g41) & (!g28) & (!g70)) + ((!g11) & (g41) & (!g28) & (g70)) + ((!g11) & (g41) & (g28) & (!g70)) + ((!g11) & (g41) & (g28) & (g70)) + ((g11) & (!g41) & (g28) & (g70)) + ((g11) & (g41) & (g28) & (g70)));
	assign g371 = (((!g25) & (!g159) & (!g368) & (!g369) & (!g370)) + ((g25) & (!g159) & (!g368) & (!g369) & (!g370)) + ((g25) & (g159) & (!g368) & (!g369) & (!g370)));
	assign g376 = (((!g50) & (g35) & (!g1) & (!g12) & (g184)) + ((!g50) & (g35) & (!g1) & (g12) & (g184)) + ((!g50) & (g35) & (g1) & (!g12) & (g184)) + ((!g50) & (g35) & (g1) & (g12) & (g184)) + ((g50) & (!g35) & (!g1) & (g12) & (!g184)) + ((g50) & (!g35) & (!g1) & (g12) & (g184)) + ((g50) & (g35) & (!g1) & (!g12) & (g184)) + ((g50) & (g35) & (!g1) & (g12) & (!g184)) + ((g50) & (g35) & (!g1) & (g12) & (g184)) + ((g50) & (g35) & (g1) & (!g12) & (g184)) + ((g50) & (g35) & (g1) & (g12) & (g184)));
	assign g381 = (((g228) & (g330) & (g371) & (g375) & (g378) & (g380)));
	assign g383 = (((!g27) & (!g45) & (!g6) & (g251) & (g287) & (!g382)) + ((!g27) & (g45) & (!g6) & (g251) & (g287) & (!g382)) + ((!g27) & (g45) & (g6) & (g251) & (g287) & (!g382)) + ((g27) & (!g45) & (!g6) & (g251) & (g287) & (!g382)) + ((g27) & (!g45) & (g6) & (g251) & (g287) & (!g382)) + ((g27) & (g45) & (!g6) & (g251) & (g287) & (!g382)) + ((g27) & (g45) & (g6) & (g251) & (g287) & (!g382)));
	assign g384 = (((!g27) & (!g42) & (g12) & (!g48) & (!g59) & (!g38)) + ((!g27) & (!g42) & (g12) & (!g48) & (!g59) & (g38)) + ((!g27) & (!g42) & (g12) & (g48) & (!g59) & (!g38)) + ((!g27) & (!g42) & (g12) & (g48) & (!g59) & (g38)) + ((!g27) & (g42) & (!g12) & (g48) & (!g59) & (!g38)) + ((!g27) & (g42) & (!g12) & (g48) & (g59) & (!g38)) + ((!g27) & (g42) & (g12) & (!g48) & (!g59) & (!g38)) + ((!g27) & (g42) & (g12) & (!g48) & (!g59) & (g38)) + ((!g27) & (g42) & (g12) & (g48) & (!g59) & (!g38)) + ((!g27) & (g42) & (g12) & (g48) & (!g59) & (g38)) + ((!g27) & (g42) & (g12) & (g48) & (g59) & (!g38)) + ((g27) & (g42) & (!g12) & (g48) & (!g59) & (!g38)) + ((g27) & (g42) & (!g12) & (g48) & (g59) & (!g38)) + ((g27) & (g42) & (g12) & (g48) & (!g59) & (!g38)) + ((g27) & (g42) & (g12) & (g48) & (g59) & (!g38)));
	assign g386 = (((!g45) & (!g1) & (!g2) & (!g38) & (!g384) & (!g385)) + ((!g45) & (!g1) & (!g2) & (g38) & (!g384) & (!g385)) + ((!g45) & (g1) & (!g2) & (!g38) & (!g384) & (!g385)) + ((!g45) & (g1) & (!g2) & (g38) & (!g384) & (!g385)) + ((!g45) & (g1) & (g2) & (!g38) & (!g384) & (!g385)) + ((!g45) & (g1) & (g2) & (g38) & (!g384) & (!g385)) + ((g45) & (!g1) & (!g2) & (!g38) & (!g384) & (!g385)) + ((g45) & (!g1) & (!g2) & (g38) & (!g384) & (!g385)) + ((g45) & (!g1) & (g2) & (g38) & (!g384) & (!g385)) + ((g45) & (g1) & (!g2) & (!g38) & (!g384) & (!g385)) + ((g45) & (g1) & (!g2) & (g38) & (!g384) & (!g385)) + ((g45) & (g1) & (g2) & (!g38) & (!g384) & (!g385)) + ((g45) & (g1) & (g2) & (g38) & (!g384) & (!g385)));
	assign g387 = (((g63) & (g42) & (g134)));
	assign g389 = (((!g28) & (!g110) & (g116) & (g141)) + ((!g28) & (g110) & (g116) & (g141)) + ((g28) & (!g110) & (g116) & (g141)) + ((g28) & (g110) & (g116) & (!g141)) + ((g28) & (g110) & (g116) & (g141)));
	assign g396 = (((!g8) & (g32) & (!g99) & (g265)) + ((!g8) & (g32) & (g99) & (g265)) + ((g8) & (!g32) & (g99) & (!g265)) + ((g8) & (!g32) & (g99) & (g265)) + ((g8) & (g32) & (!g99) & (g265)) + ((g8) & (g32) & (g99) & (!g265)) + ((g8) & (g32) & (g99) & (g265)));
	assign g398 = (((!i_3_) & (!i_5_) & (!g396) & (!g397)) + ((!i_3_) & (!i_5_) & (!g396) & (g397)) + ((!i_3_) & (i_5_) & (!g396) & (!g397)) + ((!i_3_) & (i_5_) & (!g396) & (g397)) + ((i_3_) & (!i_5_) & (!g396) & (!g397)) + ((i_3_) & (i_5_) & (!g396) & (!g397)) + ((i_3_) & (i_5_) & (!g396) & (g397)));
	assign g400 = (((!g2) & (!g3) & (!g9) & (!g243) & (g399)) + ((!g2) & (!g3) & (!g9) & (g243) & (g399)) + ((!g2) & (!g3) & (g9) & (!g243) & (g399)) + ((!g2) & (!g3) & (g9) & (g243) & (g399)) + ((!g2) & (g3) & (!g9) & (!g243) & (g399)) + ((!g2) & (g3) & (!g9) & (g243) & (g399)) + ((g2) & (!g3) & (!g9) & (!g243) & (g399)) + ((g2) & (!g3) & (g9) & (!g243) & (g399)) + ((g2) & (g3) & (!g9) & (!g243) & (g399)));
	assign g402 = (((!i_6_) & (!g25) & (g137) & (!g38) & (g401)) + ((!i_6_) & (!g25) & (g137) & (g38) & (g401)) + ((!i_6_) & (g25) & (g137) & (!g38) & (g401)) + ((!i_6_) & (g25) & (g137) & (g38) & (g401)) + ((i_6_) & (!g25) & (g137) & (!g38) & (!g401)) + ((i_6_) & (!g25) & (g137) & (!g38) & (g401)) + ((i_6_) & (!g25) & (g137) & (g38) & (g401)) + ((i_6_) & (g25) & (g137) & (!g38) & (g401)) + ((i_6_) & (g25) & (g137) & (g38) & (g401)));
	assign g405 = (((!g149) & (g398) & (g242) & (g400) & (g404)));
	assign g406 = (((i_3_) & (!i_0_) & (i_2_) & (g85)));
	assign g408 = (((!g14) & (!g1) & (!g22) & (!g406) & (!g407)) + ((!g14) & (!g1) & (!g22) & (g406) & (!g407)) + ((!g14) & (g1) & (!g22) & (!g406) & (!g407)) + ((!g14) & (g1) & (!g22) & (g406) & (!g407)) + ((!g14) & (g1) & (g22) & (!g406) & (!g407)) + ((!g14) & (g1) & (g22) & (g406) & (!g407)) + ((g14) & (!g1) & (!g22) & (!g406) & (!g407)) + ((g14) & (g1) & (!g22) & (!g406) & (!g407)) + ((g14) & (g1) & (g22) & (!g406) & (!g407)));
	assign g409 = (((!i_6_) & (!i_7_) & (i_8_) & (!g33) & (!g184) & (g401)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g33) & (g184) & (g401)) + ((!i_6_) & (!i_7_) & (i_8_) & (g33) & (!g184) & (g401)) + ((!i_6_) & (!i_7_) & (i_8_) & (g33) & (g184) & (g401)) + ((i_6_) & (!i_7_) & (i_8_) & (!g33) & (!g184) & (g401)) + ((i_6_) & (!i_7_) & (i_8_) & (!g33) & (g184) & (g401)) + ((i_6_) & (!i_7_) & (i_8_) & (g33) & (!g184) & (g401)) + ((i_6_) & (!i_7_) & (i_8_) & (g33) & (g184) & (g401)) + ((i_6_) & (i_7_) & (!i_8_) & (g33) & (!g184) & (!g401)) + ((i_6_) & (i_7_) & (!i_8_) & (g33) & (!g184) & (g401)) + ((i_6_) & (i_7_) & (!i_8_) & (g33) & (g184) & (!g401)) + ((i_6_) & (i_7_) & (!i_8_) & (g33) & (g184) & (g401)) + ((i_6_) & (i_7_) & (i_8_) & (!g33) & (g184) & (!g401)) + ((i_6_) & (i_7_) & (i_8_) & (!g33) & (g184) & (g401)) + ((i_6_) & (i_7_) & (i_8_) & (g33) & (g184) & (!g401)) + ((i_6_) & (i_7_) & (i_8_) & (g33) & (g184) & (g401)));
	assign g413 = (((g2) & (!g70) & (g158)) + ((g2) & (g70) & (!g158)) + ((g2) & (g70) & (g158)));
	assign g419 = (((!i_6_) & (!i_7_) & (i_8_) & (g189) & (!g406)) + ((!i_6_) & (!i_7_) & (i_8_) & (g189) & (g406)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g189) & (g406)) + ((!i_6_) & (i_7_) & (!i_8_) & (g189) & (g406)) + ((!i_6_) & (i_7_) & (i_8_) & (g189) & (!g406)) + ((!i_6_) & (i_7_) & (i_8_) & (g189) & (g406)) + ((i_6_) & (i_7_) & (!i_8_) & (!g189) & (g406)) + ((i_6_) & (i_7_) & (!i_8_) & (g189) & (g406)));
	assign g424 = (((!g2) & (!g38) & (!g110) & (!g421) & (g423)) + ((!g2) & (!g38) & (g110) & (!g421) & (g423)) + ((!g2) & (g38) & (!g110) & (!g421) & (g423)) + ((!g2) & (g38) & (g110) & (!g421) & (g423)) + ((g2) & (!g38) & (!g110) & (!g421) & (g423)) + ((g2) & (g38) & (!g110) & (!g421) & (g423)) + ((g2) & (g38) & (g110) & (!g421) & (g423)));
	assign g427 = (((!g24) & (!g4) & (!g425) & (!g426)) + ((g24) & (!g4) & (!g425) & (!g426)) + ((g24) & (g4) & (!g425) & (!g426)));
	assign g428 = (((!i_3_) & (i_0_) & (i_2_) & (g123)));
	assign g431 = (((!g35) & (!g1) & (g16) & (!g161)) + ((!g35) & (!g1) & (g16) & (g161)) + ((g35) & (!g1) & (!g16) & (g161)) + ((g35) & (!g1) & (g16) & (!g161)) + ((g35) & (!g1) & (g16) & (g161)) + ((g35) & (g1) & (!g16) & (g161)) + ((g35) & (g1) & (g16) & (g161)));
	assign g438 = (((!g48) & (!g33) & (!g368)) + ((!g48) & (g33) & (!g368)) + ((g48) & (!g33) & (!g368)));
	assign g445 = (((!g266) & (g438) & (g358) & (g443) & (g444)));
	assign g456 = (((!g23) & (!g66) & (!g189) & (!g455) & (!g315)) + ((g23) & (!g66) & (!g189) & (!g455) & (!g315)) + ((g23) & (!g66) & (g189) & (!g455) & (!g315)));
	assign g457 = (((!g2) & (!g36) & (!g38) & (!g110) & (g121)) + ((!g2) & (!g36) & (!g38) & (g110) & (g121)) + ((!g2) & (g36) & (!g38) & (!g110) & (g121)) + ((!g2) & (g36) & (!g38) & (g110) & (g121)) + ((g2) & (!g36) & (!g38) & (!g110) & (g121)) + ((g2) & (!g36) & (!g38) & (g110) & (!g121)) + ((g2) & (!g36) & (!g38) & (g110) & (g121)) + ((g2) & (!g36) & (g38) & (g110) & (!g121)) + ((g2) & (!g36) & (g38) & (g110) & (g121)) + ((g2) & (g36) & (!g38) & (!g110) & (g121)) + ((g2) & (g36) & (!g38) & (g110) & (g121)));
	assign g458 = (((g63) & (g64) & (g17)));
	assign g473 = (((!i_4_) & (!i_6_) & (!g4) & (!g110) & (g472)) + ((!i_4_) & (!i_6_) & (!g4) & (g110) & (g472)) + ((!i_4_) & (!i_6_) & (g4) & (!g110) & (g472)) + ((!i_4_) & (!i_6_) & (g4) & (g110) & (!g472)) + ((!i_4_) & (!i_6_) & (g4) & (g110) & (g472)) + ((!i_4_) & (i_6_) & (g4) & (g110) & (!g472)) + ((!i_4_) & (i_6_) & (g4) & (g110) & (g472)) + ((i_4_) & (!i_6_) & (g4) & (g110) & (!g472)) + ((i_4_) & (!i_6_) & (g4) & (g110) & (g472)) + ((i_4_) & (i_6_) & (g4) & (g110) & (!g472)) + ((i_4_) & (i_6_) & (g4) & (g110) & (g472)));
	assign g476 = (((!g36) & (!g121) & (g468) & (g471) & (g475)) + ((g36) & (!g121) & (g468) & (g471) & (g475)) + ((g36) & (g121) & (g468) & (g471) & (g475)));
	assign g482 = (((!g101) & (g152) & (g424) & (g480) & (g481)));
	assign g487 = (((!g155) & (!g483) & (!g484) & (!g485) & (!g486)));
	assign g491 = (((!i_5_) & (g48) & (g472)));
	assign g496 = (((!g23) & (!g91) & (!g296) & (!g491) & (g495)) + ((g23) & (!g91) & (!g296) & (!g491) & (g495)) + ((g23) & (g91) & (!g296) & (!g491) & (g495)));
	assign g497 = (((!g11) & (!i_6_) & (g2) & (!g32) & (g110)) + ((!g11) & (!i_6_) & (g2) & (g32) & (g110)) + ((!g11) & (i_6_) & (!g2) & (g32) & (g110)) + ((!g11) & (i_6_) & (g2) & (!g32) & (g110)) + ((!g11) & (i_6_) & (g2) & (g32) & (g110)) + ((g11) & (i_6_) & (!g2) & (g32) & (g110)) + ((g11) & (i_6_) & (g2) & (g32) & (g110)));
	assign g498 = (((!g35) & (!g74) & (!g189) & (!g359) & (!g497)) + ((!g35) & (!g74) & (!g189) & (g359) & (!g497)) + ((!g35) & (!g74) & (g189) & (!g359) & (!g497)) + ((!g35) & (!g74) & (g189) & (g359) & (!g497)) + ((g35) & (!g74) & (!g189) & (!g359) & (!g497)));
	assign g500 = (((!g35) & (!g25) & (!g22) & (!g36) & (!g499)) + ((!g35) & (!g25) & (!g22) & (g36) & (!g499)) + ((!g35) & (g25) & (!g22) & (!g36) & (!g499)) + ((!g35) & (g25) & (!g22) & (g36) & (!g499)) + ((!g35) & (g25) & (g22) & (!g36) & (!g499)) + ((!g35) & (g25) & (g22) & (g36) & (!g499)) + ((g35) & (!g25) & (!g22) & (g36) & (!g499)) + ((g35) & (g25) & (!g22) & (!g36) & (!g499)) + ((g35) & (g25) & (!g22) & (g36) & (!g499)) + ((g35) & (g25) & (g22) & (!g36) & (!g499)) + ((g35) & (g25) & (g22) & (g36) & (!g499)));
	assign g506 = (((!g179) & (g438) & (g498) & (g503) & (g505)));
	assign g518 = (((!g122) & (!g511) & (g513) & (g543) & (g517)));
	assign g524 = (((!g28) & (!g25) & (!g38) & (g110) & (g159)) + ((!g28) & (!g25) & (g38) & (g110) & (g159)) + ((!g28) & (g25) & (!g38) & (g110) & (g159)) + ((!g28) & (g25) & (g38) & (g110) & (g159)) + ((g28) & (!g25) & (!g38) & (!g110) & (!g159)) + ((g28) & (!g25) & (!g38) & (!g110) & (g159)) + ((g28) & (!g25) & (!g38) & (g110) & (!g159)) + ((g28) & (!g25) & (!g38) & (g110) & (g159)) + ((g28) & (!g25) & (g38) & (g110) & (g159)) + ((g28) & (g25) & (!g38) & (g110) & (g159)) + ((g28) & (g25) & (g38) & (g110) & (g159)));
	assign g528 = (((g500) & (!g525) & (!g526) & (!g527)));
	assign g531 = (((!g473) & (g498) & (!g529) & (g530)));
	assign g533 = (((!g35) & (!g23) & (!g36) & (!g110) & (g99)) + ((!g35) & (!g23) & (!g36) & (g110) & (g99)) + ((!g35) & (!g23) & (g36) & (!g110) & (g99)) + ((!g35) & (!g23) & (g36) & (g110) & (g99)) + ((g35) & (!g23) & (!g36) & (!g110) & (g99)) + ((g35) & (!g23) & (!g36) & (g110) & (!g99)) + ((g35) & (!g23) & (!g36) & (g110) & (g99)) + ((g35) & (!g23) & (g36) & (!g110) & (g99)) + ((g35) & (!g23) & (g36) & (g110) & (g99)) + ((g35) & (g23) & (!g36) & (g110) & (!g99)) + ((g35) & (g23) & (!g36) & (g110) & (g99)));
	assign g536 = (((!g28) & (!g38) & (!g110) & (!g534) & (!g535)) + ((!g28) & (!g38) & (g110) & (!g534) & (!g535)) + ((!g28) & (g38) & (!g110) & (!g534) & (!g535)) + ((!g28) & (g38) & (g110) & (!g534) & (!g535)) + ((g28) & (!g38) & (!g110) & (!g534) & (!g535)) + ((g28) & (g38) & (!g110) & (!g534) & (!g535)) + ((g28) & (g38) & (g110) & (!g534) & (!g535)));
	assign g538 = (((!g8) & (!g46) & (g2) & (g26)) + ((!g8) & (g46) & (g2) & (g26)) + ((g8) & (!g46) & (g2) & (g26)) + ((g8) & (g46) & (!g2) & (!g26)) + ((g8) & (g46) & (!g2) & (g26)) + ((g8) & (g46) & (g2) & (!g26)) + ((g8) & (g46) & (g2) & (g26)));
	assign g618 = (((!g619) & (g620)) + ((g619) & (!g620)) + ((g619) & (g620)));
	assign g631 = (((!g632) & (g633)) + ((g632) & (!g633)) + ((g632) & (g633)));
	assign g670 = (((!g671) & (g672)) + ((g671) & (!g672)) + ((g671) & (g672)));
	assign g694 = (((!g695) & (g696)) + ((g695) & (!g696)) + ((g695) & (g696)));
	assign g10 = (((!i_5_) & (g5) & (!g7) & (g9)) + ((!i_5_) & (g5) & (g7) & (g9)) + ((i_5_) & (g5) & (g7) & (!g9)) + ((i_5_) & (g5) & (g7) & (g9)));
	assign g19 = (((!g11) & (!g12) & (!g13) & (!g18)) + ((!g11) & (!g12) & (g13) & (!g18)) + ((!g11) & (g12) & (g13) & (!g18)) + ((g11) & (!g12) & (!g13) & (!g18)) + ((g11) & (!g12) & (g13) & (!g18)) + ((g11) & (g12) & (!g13) & (!g18)) + ((g11) & (g12) & (g13) & (!g18)));
	assign g39 = (((!g11) & (!g27) & (!g2) & (g37) & (!g38)) + ((!g11) & (!g27) & (g2) & (!g37) & (!g38)) + ((!g11) & (!g27) & (g2) & (!g37) & (g38)) + ((!g11) & (!g27) & (g2) & (g37) & (!g38)) + ((!g11) & (!g27) & (g2) & (g37) & (g38)) + ((g11) & (!g27) & (!g2) & (g37) & (!g38)) + ((g11) & (!g27) & (g2) & (g37) & (!g38)));
	assign g44 = (((!g11) & (!g41) & (!g43) & (!g3)) + ((!g11) & (!g41) & (!g43) & (g3)) + ((g11) & (!g41) & (!g43) & (!g3)) + ((g11) & (!g41) & (!g43) & (g3)) + ((g11) & (g41) & (!g43) & (!g3)));
	assign g53 = (((!g8) & (!g46) & (!g48) & (!g49) & (!g52)) + ((!g8) & (!g46) & (!g48) & (!g49) & (g52)) + ((!g8) & (!g46) & (!g48) & (g49) & (!g52)) + ((!g8) & (!g46) & (!g48) & (g49) & (g52)) + ((!g8) & (!g46) & (g48) & (!g49) & (!g52)) + ((!g8) & (g46) & (!g48) & (!g49) & (!g52)) + ((!g8) & (g46) & (!g48) & (!g49) & (g52)) + ((!g8) & (g46) & (!g48) & (g49) & (!g52)) + ((!g8) & (g46) & (!g48) & (g49) & (g52)) + ((!g8) & (g46) & (g48) & (!g49) & (!g52)) + ((g8) & (!g46) & (!g48) & (!g49) & (!g52)) + ((g8) & (!g46) & (!g48) & (!g49) & (g52)) + ((g8) & (!g46) & (!g48) & (g49) & (!g52)) + ((g8) & (!g46) & (!g48) & (g49) & (g52)) + ((g8) & (!g46) & (g48) & (!g49) & (!g52)));
	assign g54 = (((!i_4_) & (!i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((!i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (i_8_)) + ((!i_4_) & (i_5_) & (i_6_) & (i_7_) & (!i_8_)) + ((i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (!i_8_)) + ((i_4_) & (i_5_) & (!i_6_) & (i_7_) & (!i_8_)));
	assign g55 = (((!g50) & (g42) & (!g1) & (!g12) & (g22)) + ((!g50) & (g42) & (!g1) & (g12) & (g22)) + ((!g50) & (g42) & (g1) & (!g12) & (g22)) + ((!g50) & (g42) & (g1) & (g12) & (g22)) + ((g50) & (!g42) & (!g1) & (g12) & (!g22)) + ((g50) & (!g42) & (!g1) & (g12) & (g22)) + ((g50) & (g42) & (!g1) & (!g12) & (g22)) + ((g50) & (g42) & (!g1) & (g12) & (!g22)) + ((g50) & (g42) & (!g1) & (g12) & (g22)) + ((g50) & (g42) & (g1) & (!g12) & (g22)) + ((g50) & (g42) & (g1) & (g12) & (g22)));
	assign g56 = (((!i_3_) & (!g1) & (!g54) & (!g55)) + ((!i_3_) & (!g1) & (g54) & (!g55)) + ((!i_3_) & (g1) & (!g54) & (!g55)) + ((!i_3_) & (g1) & (g54) & (!g55)) + ((i_3_) & (!g1) & (!g54) & (!g55)) + ((i_3_) & (g1) & (!g54) & (!g55)) + ((i_3_) & (g1) & (g54) & (!g55)));
	assign g58 = (((i_4_) & (i_5_) & (g57) & (g6)));
	assign g61 = (((!g42) & (!g58) & (!g59) & (!g13) & (!g60)) + ((!g42) & (!g58) & (!g59) & (g13) & (!g60)) + ((!g42) & (!g58) & (!g59) & (g13) & (g60)) + ((!g42) & (!g58) & (g59) & (!g13) & (!g60)) + ((!g42) & (!g58) & (g59) & (!g13) & (g60)) + ((!g42) & (!g58) & (g59) & (g13) & (!g60)) + ((!g42) & (!g58) & (g59) & (g13) & (g60)) + ((g42) & (!g58) & (!g59) & (!g13) & (!g60)) + ((g42) & (!g58) & (!g59) & (g13) & (!g60)) + ((g42) & (!g58) & (g59) & (!g13) & (!g60)) + ((g42) & (!g58) & (g59) & (!g13) & (g60)) + ((g42) & (!g58) & (g59) & (g13) & (!g60)) + ((g42) & (!g58) & (g59) & (g13) & (g60)));
	assign g62 = (((g40) & (g44) & (g53) & (g56) & (g61)));
	assign g68 = (((!g1) & (!g23) & (!g32) & (!g36) & (!g67)) + ((!g1) & (!g23) & (!g32) & (!g36) & (g67)) + ((!g1) & (!g23) & (g32) & (!g36) & (!g67)) + ((!g1) & (!g23) & (g32) & (!g36) & (g67)) + ((!g1) & (!g23) & (g32) & (g36) & (g67)) + ((!g1) & (g23) & (g32) & (!g36) & (g67)) + ((!g1) & (g23) & (g32) & (g36) & (g67)) + ((g1) & (!g23) & (g32) & (!g36) & (g67)) + ((g1) & (!g23) & (g32) & (g36) & (g67)) + ((g1) & (g23) & (g32) & (!g36) & (g67)) + ((g1) & (g23) & (g32) & (g36) & (g67)));
	assign g76 = (((!g23) & (!g73) & (!g74) & (!g75)) + ((g23) & (!g73) & (!g74) & (!g75)) + ((g23) & (!g73) & (!g74) & (g75)) + ((g23) & (g73) & (!g74) & (!g75)) + ((g23) & (g73) & (!g74) & (g75)));
	assign g78 = (((!g28) & (g2) & (g77) & (!g33)) + ((!g28) & (g2) & (g77) & (g33)) + ((g28) & (!g2) & (!g77) & (g33)) + ((g28) & (!g2) & (g77) & (g33)) + ((g28) & (g2) & (!g77) & (g33)) + ((g28) & (g2) & (g77) & (!g33)) + ((g28) & (g2) & (g77) & (g33)));
	assign g79 = (((!g6) & (!g70) & (!g72) & (g76) & (!g78)) + ((!g6) & (g70) & (!g72) & (g76) & (!g78)) + ((g6) & (!g70) & (!g72) & (g76) & (!g78)));
	assign g81 = (((!g63) & (!g65) & (!g66) & (g80)) + ((!g63) & (g65) & (!g66) & (g80)) + ((g63) & (!g65) & (!g66) & (g80)));
	assign g82 = (((g20) & (g31) & (!g34) & (g62) & (g81)));
	assign g89 = (((!g23) & (!g3) & (!g29) & (g88)) + ((!g23) & (!g3) & (g29) & (g88)) + ((!g23) & (g3) & (!g29) & (g88)) + ((!g23) & (g3) & (g29) & (!g88)) + ((!g23) & (g3) & (g29) & (g88)) + ((g23) & (g3) & (g29) & (!g88)) + ((g23) & (g3) & (g29) & (g88)));
	assign g103 = (((g28) & (!g42) & (!g45) & (!g24)) + ((g28) & (g42) & (!g45) & (!g24)) + ((g28) & (g42) & (!g45) & (g24)));
	assign g104 = (((!g21) & (!g25) & (!g12) & (!g103)) + ((!g21) & (g25) & (!g12) & (!g103)) + ((!g21) & (g25) & (g12) & (!g103)) + ((g21) & (!g25) & (!g12) & (!g103)) + ((g21) & (!g25) & (g12) & (!g103)) + ((g21) & (g25) & (!g12) & (!g103)) + ((g21) & (g25) & (g12) & (!g103)));
	assign g106 = (((!g21) & (!g25) & (g48) & (!g105)) + ((!g21) & (!g25) & (g48) & (g105)) + ((!g21) & (g25) & (g48) & (!g105)) + ((g21) & (!g25) & (g48) & (!g105)) + ((g21) & (g25) & (g48) & (!g105)));
	assign g107 = (((!g35) & (!g98) & (!g102) & (g104) & (!g106)) + ((!g35) & (g98) & (!g102) & (g104) & (!g106)) + ((g35) & (!g98) & (!g102) & (g104) & (!g106)));
	assign g108 = (((!g96) & (!g97) & (!g101) & (g107)));
	assign g112 = (((!g36) & (g110) & (g111)));
	assign g113 = (((!i_7_) & (!i_8_) & (!g21) & (!g36)) + ((!i_7_) & (!i_8_) & (g21) & (!g36)) + ((i_7_) & (!i_8_) & (!g21) & (!g36)) + ((i_7_) & (!i_8_) & (!g21) & (g36)));
	assign g114 = (((!g5) & (!g36) & (!g110) & (!g111) & (!g113)) + ((!g5) & (!g36) & (!g110) & (g111) & (!g113)) + ((!g5) & (!g36) & (g110) & (!g111) & (!g113)) + ((!g5) & (g36) & (!g110) & (!g111) & (!g113)) + ((!g5) & (g36) & (!g110) & (g111) & (!g113)) + ((!g5) & (g36) & (g110) & (!g111) & (!g113)) + ((!g5) & (g36) & (g110) & (g111) & (!g113)) + ((g5) & (!g36) & (!g110) & (!g111) & (!g113)) + ((g5) & (!g36) & (g110) & (!g111) & (!g113)) + ((g5) & (g36) & (!g110) & (!g111) & (!g113)) + ((g5) & (g36) & (g110) & (!g111) & (!g113)));
	assign g115 = (((!g47) & (!g13) & (!g15) & (!g26) & (!g112) & (g114)) + ((!g47) & (!g13) & (!g15) & (!g26) & (g112) & (g114)) + ((!g47) & (!g13) & (!g15) & (g26) & (!g112) & (g114)) + ((!g47) & (!g13) & (!g15) & (g26) & (g112) & (g114)) + ((!g47) & (!g13) & (g15) & (!g26) & (!g112) & (g114)) + ((!g47) & (!g13) & (g15) & (!g26) & (g112) & (g114)) + ((!g47) & (!g13) & (g15) & (g26) & (!g112) & (g114)) + ((!g47) & (!g13) & (g15) & (g26) & (g112) & (g114)) + ((!g47) & (g13) & (!g15) & (!g26) & (!g112) & (!g114)) + ((!g47) & (g13) & (!g15) & (!g26) & (!g112) & (g114)) + ((!g47) & (g13) & (!g15) & (!g26) & (g112) & (g114)) + ((!g47) & (g13) & (!g15) & (g26) & (!g112) & (!g114)) + ((!g47) & (g13) & (!g15) & (g26) & (!g112) & (g114)) + ((!g47) & (g13) & (!g15) & (g26) & (g112) & (g114)) + ((!g47) & (g13) & (g15) & (!g26) & (!g112) & (!g114)) + ((!g47) & (g13) & (g15) & (!g26) & (!g112) & (g114)) + ((!g47) & (g13) & (g15) & (!g26) & (g112) & (g114)) + ((!g47) & (g13) & (g15) & (g26) & (!g112) & (!g114)) + ((!g47) & (g13) & (g15) & (g26) & (!g112) & (g114)) + ((!g47) & (g13) & (g15) & (g26) & (g112) & (g114)) + ((g47) & (!g13) & (!g15) & (!g26) & (!g112) & (g114)) + ((g47) & (!g13) & (!g15) & (!g26) & (g112) & (g114)) + ((g47) & (g13) & (!g15) & (!g26) & (!g112) & (!g114)) + ((g47) & (g13) & (!g15) & (!g26) & (!g112) & (g114)) + ((g47) & (g13) & (!g15) & (!g26) & (g112) & (g114)) + ((g47) & (g13) & (g15) & (!g26) & (!g112) & (!g114)) + ((g47) & (g13) & (g15) & (!g26) & (!g112) & (g114)));
	assign g118 = (((!g21) & (g42) & (!g12) & (g2) & (!g59)) + ((!g21) & (g42) & (g12) & (!g2) & (!g59)) + ((!g21) & (g42) & (g12) & (!g2) & (g59)) + ((!g21) & (g42) & (g12) & (g2) & (!g59)) + ((!g21) & (g42) & (g12) & (g2) & (g59)) + ((g21) & (g42) & (!g12) & (g2) & (!g59)) + ((g21) & (g42) & (g12) & (g2) & (!g59)));
	assign g128 = (((i_3_) & (!i_4_) & (g127)));
	assign g130 = (((!g28) & (!g75) & (!g37) & (!g99) & (!g129)) + ((!g28) & (!g75) & (!g37) & (!g99) & (g129)) + ((!g28) & (!g75) & (!g37) & (g99) & (!g129)) + ((!g28) & (!g75) & (!g37) & (g99) & (g129)) + ((!g28) & (!g75) & (g37) & (!g99) & (!g129)) + ((!g28) & (!g75) & (g37) & (g99) & (!g129)) + ((!g28) & (g75) & (!g37) & (!g99) & (!g129)) + ((!g28) & (g75) & (!g37) & (!g99) & (g129)) + ((!g28) & (g75) & (!g37) & (g99) & (!g129)) + ((!g28) & (g75) & (!g37) & (g99) & (g129)) + ((!g28) & (g75) & (g37) & (!g99) & (!g129)) + ((!g28) & (g75) & (g37) & (g99) & (!g129)) + ((g28) & (!g75) & (!g37) & (!g99) & (!g129)) + ((g28) & (!g75) & (g37) & (!g99) & (!g129)));
	assign g131 = (((!g120) & (!g1) & (!g48) & (g2) & (!g38)) + ((!g120) & (!g1) & (g48) & (g2) & (!g38)) + ((g120) & (!g1) & (!g48) & (g2) & (!g38)) + ((g120) & (!g1) & (g48) & (!g2) & (!g38)) + ((g120) & (!g1) & (g48) & (!g2) & (g38)) + ((g120) & (!g1) & (g48) & (g2) & (!g38)) + ((g120) & (!g1) & (g48) & (g2) & (g38)));
	assign g132 = (((!g12) & (g683) & (!g128) & (g130) & (!g131)) + ((!g12) & (g683) & (g128) & (g130) & (!g131)) + ((g12) & (g683) & (!g128) & (g130) & (!g131)));
	assign g133 = (((g694) & (!g122) & (g125) & (g132)));
	assign g136 = (((!i_3_) & (!i_5_) & (!i_2_) & (g35) & (!g14) & (!g64)) + ((!i_3_) & (!i_5_) & (!i_2_) & (g35) & (!g14) & (g64)) + ((!i_3_) & (!i_5_) & (!i_2_) & (g35) & (g14) & (!g64)) + ((!i_3_) & (!i_5_) & (!i_2_) & (g35) & (g14) & (g64)) + ((i_3_) & (!i_5_) & (i_2_) & (!g35) & (g14) & (g64)) + ((i_3_) & (!i_5_) & (i_2_) & (g35) & (g14) & (g64)) + ((i_3_) & (i_5_) & (i_2_) & (!g35) & (g14) & (g64)) + ((i_3_) & (i_5_) & (i_2_) & (g35) & (g14) & (g64)));
	assign g138 = (((!i_3_) & (!i_0_) & (i_1_) & (g137) & (g85)));
	assign g139 = (((!i_3_) & (i_5_) & (g28) & (!g24)));
	assign g142 = (((!i_3_) & (!g42) & (!g8) & (!g45) & (g141)) + ((!i_3_) & (!g42) & (g8) & (!g45) & (g141)) + ((!i_3_) & (g42) & (!g8) & (!g45) & (g141)) + ((!i_3_) & (g42) & (g8) & (!g45) & (!g141)) + ((!i_3_) & (g42) & (g8) & (!g45) & (g141)) + ((!i_3_) & (g42) & (g8) & (g45) & (!g141)) + ((!i_3_) & (g42) & (g8) & (g45) & (g141)) + ((i_3_) & (!g42) & (!g8) & (!g45) & (g141)) + ((i_3_) & (!g42) & (g8) & (!g45) & (g141)) + ((i_3_) & (g42) & (!g8) & (!g45) & (g141)) + ((i_3_) & (g42) & (g8) & (!g45) & (g141)));
	assign g143 = (((!i_8_) & (!g51) & (!g64) & (!g142)) + ((!i_8_) & (!g51) & (g64) & (!g142)) + ((!i_8_) & (g51) & (!g64) & (!g142)) + ((i_8_) & (!g51) & (!g64) & (!g142)) + ((i_8_) & (!g51) & (g64) & (!g142)) + ((i_8_) & (g51) & (!g64) & (!g142)) + ((i_8_) & (g51) & (g64) & (!g142)));
	assign g144 = (((!i_1_) & (!g135) & (!g136) & (g140) & (g143)) + ((!i_1_) & (!g135) & (g136) & (g140) & (g143)) + ((!i_1_) & (g135) & (!g136) & (g140) & (g143)) + ((!i_1_) & (g135) & (g136) & (g140) & (g143)) + ((i_1_) & (!g135) & (!g136) & (g140) & (g143)));
	assign g146 = (((!g27) & (!i_6_) & (g47) & (!g24) & (g3)) + ((!g27) & (!i_6_) & (g47) & (g24) & (g3)) + ((!g27) & (i_6_) & (g47) & (!g24) & (g3)) + ((!g27) & (i_6_) & (g47) & (g24) & (g3)) + ((g27) & (i_6_) & (g47) & (!g24) & (g3)));
	assign g148 = (((!g11) & (g42) & (!g47) & (!g64) & (g111)) + ((!g11) & (g42) & (!g47) & (g64) & (g111)) + ((!g11) & (g42) & (g47) & (!g64) & (g111)) + ((!g11) & (g42) & (g47) & (g64) & (!g111)) + ((!g11) & (g42) & (g47) & (g64) & (g111)) + ((g11) & (g42) & (g47) & (g64) & (!g111)) + ((g11) & (g42) & (g47) & (g64) & (g111)));
	assign g151 = (((!g25) & (!g12) & (!g3) & (!g150)) + ((!g25) & (!g12) & (g3) & (!g150)) + ((!g25) & (g12) & (!g3) & (!g150)) + ((g25) & (!g12) & (!g3) & (!g150)) + ((g25) & (!g12) & (g3) & (!g150)) + ((g25) & (g12) & (!g3) & (!g150)) + ((g25) & (g12) & (g3) & (!g150)));
	assign g153 = (((g670) & (g147) & (g152)));
	assign g156 = (((!g23) & (!g36) & (!g7) & (g129)) + ((!g23) & (!g36) & (g7) & (!g129)) + ((!g23) & (!g36) & (g7) & (g129)) + ((!g23) & (g36) & (!g7) & (g129)) + ((!g23) & (g36) & (g7) & (g129)) + ((g23) & (!g36) & (g7) & (!g129)) + ((g23) & (!g36) & (g7) & (g129)));
	assign g162 = (((!g28) & (g2) & (!g24) & (g32) & (!g161)) + ((!g28) & (g2) & (!g24) & (g32) & (g161)) + ((g28) & (!g2) & (!g24) & (!g32) & (g161)) + ((g28) & (!g2) & (!g24) & (g32) & (g161)) + ((g28) & (!g2) & (g24) & (!g32) & (g161)) + ((g28) & (!g2) & (g24) & (g32) & (g161)) + ((g28) & (g2) & (!g24) & (!g32) & (g161)) + ((g28) & (g2) & (!g24) & (g32) & (!g161)) + ((g28) & (g2) & (!g24) & (g32) & (g161)) + ((g28) & (g2) & (g24) & (!g32) & (g161)) + ((g28) & (g2) & (g24) & (g32) & (g161)));
	assign g163 = (((i_7_) & (!i_8_) & (!g45) & (!g13) & (!g88)) + ((i_7_) & (!i_8_) & (!g45) & (!g13) & (g88)) + ((i_7_) & (i_8_) & (!g45) & (!g13) & (g88)) + ((i_7_) & (i_8_) & (!g45) & (g13) & (g88)) + ((i_7_) & (i_8_) & (g45) & (!g13) & (g88)) + ((i_7_) & (i_8_) & (g45) & (g13) & (g88)));
	assign g169 = (((g50) & (i_6_) & (g42) & (g47)));
	assign g171 = (((!i_3_) & (i_5_) & (g2) & (!g13)));
	assign g172 = (((!g32) & (!g121) & (!g170) & (!g171)) + ((!g32) & (g121) & (!g170) & (!g171)) + ((g32) & (!g121) & (!g170) & (!g171)));
	assign g176 = (((!g28) & (!g25) & (!g59) & (g7) & (!g110)) + ((!g28) & (!g25) & (!g59) & (g7) & (g110)) + ((!g28) & (g25) & (!g59) & (g7) & (!g110)) + ((!g28) & (g25) & (!g59) & (g7) & (g110)) + ((g28) & (!g25) & (!g59) & (!g7) & (!g110)) + ((g28) & (!g25) & (!g59) & (!g7) & (g110)) + ((g28) & (!g25) & (!g59) & (g7) & (!g110)) + ((g28) & (!g25) & (!g59) & (g7) & (g110)) + ((g28) & (g25) & (!g59) & (!g7) & (g110)) + ((g28) & (g25) & (!g59) & (g7) & (!g110)) + ((g28) & (g25) & (!g59) & (g7) & (g110)));
	assign g177 = (((!g173) & (!g174) & (!g175) & (!g176)));
	assign g180 = (((!i_3_) & (!i_4_) & (i_5_) & (!g127) & (g63) & (g51)) + ((!i_3_) & (!i_4_) & (i_5_) & (g127) & (g63) & (g51)) + ((i_3_) & (!i_4_) & (i_5_) & (!g127) & (g63) & (g51)) + ((i_3_) & (!i_4_) & (i_5_) & (g127) & (g63) & (g51)) + ((i_3_) & (i_4_) & (i_5_) & (g127) & (g63) & (!g51)) + ((i_3_) & (i_4_) & (i_5_) & (g127) & (g63) & (g51)));
	assign g182 = (((!i_6_) & (i_7_) & (!i_8_) & (g75) & (!g181) & (!g105)) + ((!i_6_) & (i_7_) & (!i_8_) & (g75) & (!g181) & (g105)) + ((!i_6_) & (i_7_) & (!i_8_) & (g75) & (g181) & (!g105)) + ((!i_6_) & (i_7_) & (!i_8_) & (g75) & (g181) & (g105)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g75) & (!g181) & (!g105)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g75) & (g181) & (!g105)) + ((i_6_) & (!i_7_) & (!i_8_) & (g75) & (!g181) & (!g105)) + ((i_6_) & (!i_7_) & (!i_8_) & (g75) & (g181) & (!g105)) + ((i_6_) & (i_7_) & (i_8_) & (!g75) & (g181) & (!g105)) + ((i_6_) & (i_7_) & (i_8_) & (!g75) & (g181) & (g105)) + ((i_6_) & (i_7_) & (i_8_) & (g75) & (g181) & (!g105)) + ((i_6_) & (i_7_) & (i_8_) & (g75) & (g181) & (g105)));
	assign g183 = (((!i_3_) & (!i_5_) & (g127) & (!g28) & (g123)) + ((!i_3_) & (!i_5_) & (g127) & (g28) & (g123)) + ((!i_3_) & (i_5_) & (g127) & (!g28) & (g123)) + ((!i_3_) & (i_5_) & (g127) & (g28) & (g123)) + ((i_3_) & (i_5_) & (g127) & (g28) & (!g123)) + ((i_3_) & (i_5_) & (g127) & (g28) & (g123)));
	assign g185 = (((!g2) & (!g23) & (!g70) & (g184)) + ((!g2) & (!g23) & (g70) & (g184)) + ((g2) & (!g23) & (!g70) & (g184)) + ((g2) & (!g23) & (g70) & (!g184)) + ((g2) & (!g23) & (g70) & (g184)) + ((g2) & (g23) & (g70) & (!g184)) + ((g2) & (g23) & (g70) & (g184)));
	assign g190 = (((!i_6_) & (!g63) & (!g188) & (!g181) & (!g189)) + ((!i_6_) & (!g63) & (!g188) & (!g181) & (g189)) + ((!i_6_) & (!g63) & (!g188) & (g181) & (!g189)) + ((!i_6_) & (!g63) & (!g188) & (g181) & (g189)) + ((!i_6_) & (g63) & (!g188) & (!g181) & (!g189)) + ((!i_6_) & (g63) & (!g188) & (g181) & (!g189)) + ((i_6_) & (!g63) & (!g188) & (!g181) & (!g189)) + ((i_6_) & (!g63) & (!g188) & (!g181) & (g189)) + ((i_6_) & (!g63) & (!g188) & (g181) & (!g189)) + ((i_6_) & (!g63) & (!g188) & (g181) & (g189)) + ((i_6_) & (g63) & (!g188) & (!g181) & (!g189)) + ((i_6_) & (g63) & (!g188) & (!g181) & (g189)));
	assign g191 = (((!g185) & (!g186) & (g657) & (g190)));
	assign g192 = (((!g179) & (!g180) & (!g182) & (!g183) & (g191)));
	assign g196 = (((!g27) & (!g23) & (!g3) & (g110) & (g194)) + ((!g27) & (!g23) & (g3) & (!g110) & (!g194)) + ((!g27) & (!g23) & (g3) & (!g110) & (g194)) + ((!g27) & (!g23) & (g3) & (g110) & (!g194)) + ((!g27) & (!g23) & (g3) & (g110) & (g194)) + ((!g27) & (g23) & (!g3) & (g110) & (g194)) + ((!g27) & (g23) & (g3) & (g110) & (g194)) + ((g27) & (!g23) & (!g3) & (g110) & (g194)) + ((g27) & (!g23) & (g3) & (g110) & (g194)) + ((g27) & (g23) & (!g3) & (g110) & (g194)) + ((g27) & (g23) & (g3) & (g110) & (g194)));
	assign g197 = (((!g47) & (!g73) & (!g193) & (!g195) & (!g196)) + ((!g47) & (g73) & (!g193) & (!g195) & (!g196)) + ((g47) & (!g73) & (!g193) & (!g195) & (!g196)));
	assign g198 = (((g166) & (!g168) & (g178) & (g192) & (g197)));
	assign g199 = (((g109) & (g154) & (g157) & (g164) & (g198)));
	assign g201 = (((!g50) & (!i_6_) & (g137) & (!g94) & (g88)) + ((!g50) & (!i_6_) & (g137) & (g94) & (g88)) + ((g50) & (!i_6_) & (g137) & (!g94) & (g88)) + ((g50) & (!i_6_) & (g137) & (g94) & (g88)) + ((g50) & (i_6_) & (g137) & (g94) & (!g88)) + ((g50) & (i_6_) & (g137) & (g94) & (g88)));
	assign g203 = (((!i_6_) & (g63) & (!g21) & (!g13) & (!g84)) + ((!i_6_) & (g63) & (!g21) & (!g13) & (g84)) + ((i_6_) & (g63) & (!g21) & (!g13) & (g84)) + ((i_6_) & (g63) & (!g21) & (g13) & (g84)) + ((i_6_) & (g63) & (g21) & (!g13) & (g84)) + ((i_6_) & (g63) & (g21) & (g13) & (g84)));
	assign g205 = (((!g23) & (!g70) & (!g204)) + ((g23) & (!g70) & (!g204)) + ((g23) & (g70) & (!g204)));
	assign g207 = (((!i_3_) & (!i_5_) & (g8) & (!g24)));
	assign g209 = (((g127) & (!i_2_) & (!g8) & (g22) & (!g59)) + ((g127) & (!i_2_) & (!g8) & (g22) & (g59)) + ((g127) & (!i_2_) & (g8) & (g22) & (!g59)) + ((g127) & (!i_2_) & (g8) & (g22) & (g59)) + ((g127) & (i_2_) & (g8) & (!g22) & (!g59)) + ((g127) & (i_2_) & (g8) & (g22) & (!g59)));
	assign g210 = (((!g28) & (!g26) & (!g208) & (g644) & (!g209)) + ((!g28) & (g26) & (!g208) & (g644) & (!g209)) + ((g28) & (!g26) & (!g208) & (g644) & (!g209)));
	assign g213 = (((g50) & (i_6_) & (g42) & (g137)));
	assign g214 = (((!g2) & (!g73) & (!g38) & (!g29) & (!g213)) + ((!g2) & (!g73) & (g38) & (!g29) & (!g213)) + ((!g2) & (!g73) & (g38) & (g29) & (!g213)) + ((!g2) & (g73) & (!g38) & (!g29) & (!g213)) + ((!g2) & (g73) & (g38) & (!g29) & (!g213)) + ((!g2) & (g73) & (g38) & (g29) & (!g213)) + ((g2) & (!g73) & (!g38) & (!g29) & (!g213)) + ((g2) & (!g73) & (g38) & (!g29) & (!g213)) + ((g2) & (!g73) & (g38) & (g29) & (!g213)));
	assign g220 = (((!i_3_) & (i_1_) & (!i_2_) & (g219)));
	assign g221 = (((!g27) & (!g35) & (g28) & (!g1) & (!g36)) + ((!g27) & (!g35) & (g28) & (g1) & (!g36)) + ((!g27) & (g35) & (!g28) & (!g1) & (!g36)) + ((!g27) & (g35) & (g28) & (!g1) & (!g36)) + ((!g27) & (g35) & (g28) & (g1) & (!g36)) + ((g27) & (g35) & (!g28) & (!g1) & (!g36)) + ((g27) & (g35) & (g28) & (!g1) & (!g36)));
	assign g222 = (((!g23) & (!g59) & (g13) & (g105) & (!g221)) + ((!g23) & (g59) & (!g13) & (g105) & (!g221)) + ((!g23) & (g59) & (g13) & (g105) & (!g221)) + ((g23) & (!g59) & (!g13) & (!g105) & (!g221)) + ((g23) & (!g59) & (!g13) & (g105) & (!g221)) + ((g23) & (!g59) & (g13) & (!g105) & (!g221)) + ((g23) & (!g59) & (g13) & (g105) & (!g221)) + ((g23) & (g59) & (!g13) & (!g105) & (!g221)) + ((g23) & (g59) & (!g13) & (g105) & (!g221)) + ((g23) & (g59) & (g13) & (!g105) & (!g221)) + ((g23) & (g59) & (g13) & (g105) & (!g221)));
	assign g223 = (((!g27) & (!g43) & (!g23) & (!g3)) + ((!g27) & (!g43) & (g23) & (!g3)) + ((!g27) & (!g43) & (g23) & (g3)) + ((g27) & (!g43) & (!g23) & (!g3)) + ((g27) & (!g43) & (!g23) & (g3)) + ((g27) & (!g43) & (g23) & (!g3)) + ((g27) & (!g43) & (g23) & (g3)));
	assign g227 = (((!i_6_) & (!i_7_) & (i_8_) & (g100) & (!g129)) + ((!i_6_) & (!i_7_) & (i_8_) & (g100) & (g129)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g100) & (g129)));
	assign g231 = (((g50) & (!g8) & (g12) & (!g57) & (g230)) + ((g50) & (!g8) & (g12) & (g57) & (g230)) + ((g50) & (g8) & (!g12) & (g57) & (!g230)) + ((g50) & (g8) & (!g12) & (g57) & (g230)) + ((g50) & (g8) & (g12) & (!g57) & (g230)) + ((g50) & (g8) & (g12) & (g57) & (!g230)) + ((g50) & (g8) & (g12) & (g57) & (g230)));
	assign g232 = (((!i_6_) & (!i_7_) & (!i_8_) & (!g75) & (!g158) & (!g231)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g75) & (!g158) & (!g231)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g75) & (!g158) & (!g231)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g75) & (g158) & (!g231)) + ((!i_6_) & (!i_7_) & (i_8_) & (g75) & (!g158) & (!g231)) + ((!i_6_) & (!i_7_) & (i_8_) & (g75) & (g158) & (!g231)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g75) & (!g158) & (!g231)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g75) & (g158) & (!g231)) + ((!i_6_) & (i_7_) & (i_8_) & (!g75) & (!g158) & (!g231)) + ((!i_6_) & (i_7_) & (i_8_) & (!g75) & (g158) & (!g231)) + ((!i_6_) & (i_7_) & (i_8_) & (g75) & (!g158) & (!g231)) + ((!i_6_) & (i_7_) & (i_8_) & (g75) & (g158) & (!g231)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g75) & (!g158) & (!g231)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g75) & (g158) & (!g231)) + ((i_6_) & (!i_7_) & (i_8_) & (!g75) & (!g158) & (!g231)) + ((i_6_) & (!i_7_) & (i_8_) & (!g75) & (g158) & (!g231)) + ((i_6_) & (!i_7_) & (i_8_) & (g75) & (!g158) & (!g231)) + ((i_6_) & (!i_7_) & (i_8_) & (g75) & (g158) & (!g231)) + ((i_6_) & (i_7_) & (!i_8_) & (!g75) & (!g158) & (!g231)) + ((i_6_) & (i_7_) & (!i_8_) & (!g75) & (g158) & (!g231)) + ((i_6_) & (i_7_) & (!i_8_) & (g75) & (!g158) & (!g231)) + ((i_6_) & (i_7_) & (!i_8_) & (g75) & (g158) & (!g231)) + ((i_6_) & (i_7_) & (i_8_) & (!g75) & (!g158) & (!g231)) + ((i_6_) & (i_7_) & (i_8_) & (!g75) & (g158) & (!g231)));
	assign g233 = (((!g25) & (!g194) & (!g229) & (g631) & (g232)) + ((g25) & (!g194) & (!g229) & (g631) & (g232)) + ((g25) & (g194) & (!g229) & (g631) & (g232)));
	assign g235 = (((!g35) & (!g21) & (g8) & (!g25) & (g32)) + ((!g35) & (g21) & (g8) & (!g25) & (g32)) + ((g35) & (!g21) & (!g8) & (!g25) & (!g32)) + ((g35) & (!g21) & (!g8) & (!g25) & (g32)) + ((g35) & (!g21) & (g8) & (!g25) & (!g32)) + ((g35) & (!g21) & (g8) & (!g25) & (g32)) + ((g35) & (g21) & (g8) & (!g25) & (g32)));
	assign g237 = (((!g21) & (!g8) & (!g24) & (g69)) + ((!g21) & (!g8) & (g24) & (g69)) + ((!g21) & (g8) & (g24) & (g69)) + ((g21) & (!g8) & (!g24) & (g69)) + ((g21) & (!g8) & (g24) & (g69)) + ((g21) & (g8) & (!g24) & (g69)) + ((g21) & (g8) & (g24) & (g69)));
	assign g238 = (((!g11) & (!g1) & (!g23) & (!g3) & (g141)) + ((!g11) & (!g1) & (!g23) & (g3) & (!g141)) + ((!g11) & (!g1) & (!g23) & (g3) & (g141)) + ((!g11) & (!g1) & (g23) & (!g3) & (g141)) + ((!g11) & (!g1) & (g23) & (g3) & (g141)) + ((!g11) & (g1) & (!g23) & (!g3) & (g141)) + ((!g11) & (g1) & (!g23) & (g3) & (g141)) + ((!g11) & (g1) & (g23) & (!g3) & (g141)) + ((!g11) & (g1) & (g23) & (g3) & (g141)) + ((g11) & (!g1) & (!g23) & (g3) & (!g141)) + ((g11) & (!g1) & (!g23) & (g3) & (g141)));
	assign g240 = (((!g25) & (!g120) & (g12) & (g181)) + ((!g25) & (g120) & (g12) & (!g181)) + ((!g25) & (g120) & (g12) & (g181)) + ((g25) & (!g120) & (g12) & (g181)) + ((g25) & (g120) & (g12) & (g181)));
	assign g241 = (((!g59) & (!g29) & (!g239) & (!g240)) + ((g59) & (!g29) & (!g239) & (!g240)) + ((g59) & (g29) & (!g239) & (!g240)));
	assign g245 = (((!g2) & (!g24) & (!g32) & (!g244)) + ((!g2) & (!g24) & (g32) & (!g244)) + ((!g2) & (g24) & (!g32) & (!g244)) + ((!g2) & (g24) & (g32) & (!g244)) + ((g2) & (!g24) & (!g32) & (!g244)) + ((g2) & (g24) & (!g32) & (!g244)) + ((g2) & (g24) & (g32) & (!g244)));
	assign g248 = (((!g45) & (!g38) & (!g29) & (g121)) + ((!g45) & (!g38) & (g29) & (!g121)) + ((!g45) & (!g38) & (g29) & (g121)) + ((!g45) & (g38) & (g29) & (!g121)) + ((!g45) & (g38) & (g29) & (g121)) + ((g45) & (!g38) & (!g29) & (g121)) + ((g45) & (!g38) & (g29) & (g121)));
	assign g250 = (((i_3_) & (!i_4_) & (!g27) & (i_6_) & (!i_8_)));
	assign g253 = (((!g48) & (!g57) & (!g33) & (!g16) & (!g252)) + ((!g48) & (!g57) & (!g33) & (g16) & (!g252)) + ((!g48) & (!g57) & (g33) & (!g16) & (!g252)) + ((!g48) & (!g57) & (g33) & (g16) & (!g252)) + ((!g48) & (g57) & (!g33) & (!g16) & (!g252)) + ((!g48) & (g57) & (g33) & (!g16) & (!g252)) + ((g48) & (!g57) & (!g33) & (!g16) & (!g252)) + ((g48) & (!g57) & (!g33) & (g16) & (!g252)) + ((g48) & (g57) & (!g33) & (!g16) & (!g252)));
	assign g258 = (((!g28) & (!g70) & (!g189) & (!g167) & (!g230)) + ((!g28) & (!g70) & (!g189) & (!g167) & (g230)) + ((!g28) & (!g70) & (!g189) & (g167) & (!g230)) + ((!g28) & (!g70) & (g189) & (!g167) & (!g230)) + ((!g28) & (!g70) & (g189) & (!g167) & (g230)) + ((!g28) & (!g70) & (g189) & (g167) & (!g230)) + ((!g28) & (g70) & (!g189) & (!g167) & (!g230)) + ((!g28) & (g70) & (!g189) & (!g167) & (g230)) + ((!g28) & (g70) & (!g189) & (g167) & (!g230)) + ((!g28) & (g70) & (g189) & (!g167) & (!g230)) + ((!g28) & (g70) & (g189) & (!g167) & (g230)) + ((!g28) & (g70) & (g189) & (g167) & (!g230)) + ((g28) & (!g70) & (!g189) & (!g167) & (!g230)) + ((g28) & (!g70) & (!g189) & (!g167) & (g230)) + ((g28) & (!g70) & (!g189) & (g167) & (!g230)));
	assign g259 = (((!g45) & (!g6) & (!g110) & (g141)) + ((!g45) & (!g6) & (g110) & (g141)) + ((!g45) & (g6) & (!g110) & (g141)) + ((!g45) & (g6) & (g110) & (!g141)) + ((!g45) & (g6) & (g110) & (g141)));
	assign g260 = (((!g24) & (!g36) & (!g60) & (!g4) & (!g259)) + ((!g24) & (g36) & (!g60) & (!g4) & (!g259)) + ((!g24) & (g36) & (g60) & (!g4) & (!g259)) + ((g24) & (!g36) & (!g60) & (!g4) & (!g259)) + ((g24) & (!g36) & (!g60) & (g4) & (!g259)) + ((g24) & (!g36) & (g60) & (!g4) & (!g259)) + ((g24) & (!g36) & (g60) & (g4) & (!g259)) + ((g24) & (g36) & (!g60) & (!g4) & (!g259)) + ((g24) & (g36) & (!g60) & (g4) & (!g259)) + ((g24) & (g36) & (g60) & (!g4) & (!g259)) + ((g24) & (g36) & (g60) & (g4) & (!g259)));
	assign g261 = (((!g83) & (!g255) & (g257) & (g258) & (g260)));
	assign g262 = (((g237) & (g242) & (g246) & (g249) & (g254) & (g261)));
	assign g263 = (((g157) & (g206) & (g211) & (g234) & (g236) & (g262)));
	assign g269 = (((!i_7_) & (g28) & (g75) & (!g268)) + ((!i_7_) & (g28) & (g75) & (g268)) + ((i_7_) & (!g28) & (!g75) & (g268)) + ((i_7_) & (!g28) & (g75) & (g268)) + ((i_7_) & (g28) & (!g75) & (g268)) + ((i_7_) & (g28) & (g75) & (!g268)) + ((i_7_) & (g28) & (g75) & (g268)));
	assign g270 = (((!g1) & (g6) & (!g36) & (!g49)) + ((!g1) & (g6) & (!g36) & (g49)) + ((!g1) & (g6) & (g36) & (g49)) + ((g1) & (g6) & (!g36) & (g49)) + ((g1) & (g6) & (g36) & (g49)));
	assign g271 = (((!g27) & (!g45) & (!g1) & (!g23) & (!g4) & (!g189)) + ((!g27) & (!g45) & (!g1) & (!g23) & (!g4) & (g189)) + ((!g27) & (!g45) & (!g1) & (!g23) & (g4) & (!g189)) + ((!g27) & (!g45) & (!g1) & (!g23) & (g4) & (g189)) + ((!g27) & (!g45) & (!g1) & (g23) & (g4) & (!g189)) + ((!g27) & (!g45) & (!g1) & (g23) & (g4) & (g189)) + ((!g27) & (!g45) & (g1) & (!g23) & (!g4) & (g189)) + ((!g27) & (!g45) & (g1) & (!g23) & (g4) & (!g189)) + ((!g27) & (!g45) & (g1) & (!g23) & (g4) & (g189)) + ((!g27) & (!g45) & (g1) & (g23) & (g4) & (!g189)) + ((!g27) & (!g45) & (g1) & (g23) & (g4) & (g189)) + ((!g27) & (g45) & (!g1) & (!g23) & (!g4) & (g189)) + ((!g27) & (g45) & (!g1) & (!g23) & (g4) & (!g189)) + ((!g27) & (g45) & (!g1) & (!g23) & (g4) & (g189)) + ((!g27) & (g45) & (!g1) & (g23) & (g4) & (!g189)) + ((!g27) & (g45) & (!g1) & (g23) & (g4) & (g189)) + ((!g27) & (g45) & (g1) & (!g23) & (!g4) & (g189)) + ((!g27) & (g45) & (g1) & (!g23) & (g4) & (!g189)) + ((!g27) & (g45) & (g1) & (!g23) & (g4) & (g189)) + ((!g27) & (g45) & (g1) & (g23) & (g4) & (!g189)) + ((!g27) & (g45) & (g1) & (g23) & (g4) & (g189)) + ((g27) & (!g45) & (!g1) & (!g23) & (!g4) & (!g189)) + ((g27) & (!g45) & (!g1) & (!g23) & (!g4) & (g189)) + ((g27) & (!g45) & (!g1) & (!g23) & (g4) & (!g189)) + ((g27) & (!g45) & (!g1) & (!g23) & (g4) & (g189)) + ((g27) & (!g45) & (g1) & (!g23) & (!g4) & (g189)) + ((g27) & (!g45) & (g1) & (!g23) & (g4) & (g189)) + ((g27) & (g45) & (!g1) & (!g23) & (!g4) & (g189)) + ((g27) & (g45) & (!g1) & (!g23) & (g4) & (g189)) + ((g27) & (g45) & (g1) & (!g23) & (!g4) & (g189)) + ((g27) & (g45) & (g1) & (!g23) & (g4) & (g189)));
	assign g272 = (((!g48) & (!g105) & (!g270) & (!g271)) + ((!g48) & (g105) & (!g270) & (!g271)) + ((g48) & (g105) & (!g270) & (!g271)));
	assign g273 = (((!g8) & (!g77) & (!g200) & (!g269) & (g272)) + ((!g8) & (g77) & (!g200) & (!g269) & (g272)) + ((g8) & (!g77) & (!g200) & (!g269) & (g272)));
	assign g280 = (((!g25) & (!g6) & (!g32) & (!g121) & (!g252)) + ((!g25) & (!g6) & (!g32) & (g121) & (!g252)) + ((!g25) & (!g6) & (g32) & (!g121) & (!g252)) + ((!g25) & (g6) & (!g32) & (!g121) & (!g252)) + ((!g25) & (g6) & (!g32) & (g121) & (!g252)) + ((g25) & (!g6) & (!g32) & (!g121) & (!g252)) + ((g25) & (!g6) & (!g32) & (g121) & (!g252)) + ((g25) & (!g6) & (g32) & (!g121) & (!g252)) + ((g25) & (g6) & (!g32) & (!g121) & (!g252)) + ((g25) & (g6) & (!g32) & (g121) & (!g252)) + ((g25) & (g6) & (g32) & (!g121) & (!g252)));
	assign g281 = (((!g35) & (g6) & (!g117) & (g161)) + ((!g35) & (g6) & (g117) & (g161)) + ((g35) & (!g6) & (g117) & (!g161)) + ((g35) & (!g6) & (g117) & (g161)) + ((g35) & (g6) & (!g117) & (g161)) + ((g35) & (g6) & (g117) & (!g161)) + ((g35) & (g6) & (g117) & (g161)));
	assign g282 = (((!g277) & (!g278) & (!g279) & (g280) & (!g281)));
	assign g284 = (((!g27) & (g137) & (g15)));
	assign g286 = (((!g2) & (!g26) & (!g155)) + ((!g2) & (g26) & (!g155)) + ((g2) & (!g26) & (!g155)));
	assign g288 = (((!g28) & (g12) & (g184) & (!g243)) + ((!g28) & (g12) & (g184) & (g243)) + ((g28) & (!g12) & (!g184) & (g243)) + ((g28) & (!g12) & (g184) & (g243)) + ((g28) & (g12) & (!g184) & (g243)) + ((g28) & (g12) & (g184) & (!g243)) + ((g28) & (g12) & (g184) & (g243)));
	assign g295 = (((!i_5_) & (!g35) & (!g42) & (!g5) & (!g121) & (!g294)) + ((!i_5_) & (!g35) & (!g42) & (!g5) & (g121) & (!g294)) + ((!i_5_) & (!g35) & (!g42) & (g5) & (!g121) & (!g294)) + ((!i_5_) & (!g35) & (!g42) & (g5) & (g121) & (!g294)) + ((!i_5_) & (!g35) & (g42) & (!g5) & (!g121) & (!g294)) + ((!i_5_) & (!g35) & (g42) & (!g5) & (g121) & (!g294)) + ((!i_5_) & (!g35) & (g42) & (g5) & (!g121) & (!g294)) + ((!i_5_) & (!g35) & (g42) & (g5) & (g121) & (!g294)) + ((!i_5_) & (g35) & (!g42) & (!g5) & (!g121) & (!g294)) + ((!i_5_) & (g35) & (!g42) & (!g5) & (g121) & (!g294)) + ((!i_5_) & (g35) & (!g42) & (g5) & (!g121) & (!g294)) + ((!i_5_) & (g35) & (!g42) & (g5) & (g121) & (!g294)) + ((!i_5_) & (g35) & (g42) & (!g5) & (!g121) & (!g294)) + ((!i_5_) & (g35) & (g42) & (!g5) & (g121) & (!g294)) + ((i_5_) & (!g35) & (!g42) & (!g5) & (!g121) & (!g294)) + ((i_5_) & (!g35) & (!g42) & (!g5) & (g121) & (!g294)) + ((i_5_) & (!g35) & (!g42) & (g5) & (!g121) & (!g294)) + ((i_5_) & (!g35) & (g42) & (!g5) & (!g121) & (!g294)) + ((i_5_) & (!g35) & (g42) & (!g5) & (g121) & (!g294)) + ((i_5_) & (!g35) & (g42) & (g5) & (!g121) & (!g294)) + ((i_5_) & (g35) & (!g42) & (!g5) & (!g121) & (!g294)) + ((i_5_) & (g35) & (!g42) & (!g5) & (g121) & (!g294)) + ((i_5_) & (g35) & (!g42) & (g5) & (!g121) & (!g294)) + ((i_5_) & (g35) & (g42) & (!g5) & (!g121) & (!g294)) + ((i_5_) & (g35) & (g42) & (!g5) & (g121) & (!g294)) + ((i_5_) & (g35) & (g42) & (g5) & (!g121) & (!g294)));
	assign g297 = (((!i_3_) & (!i_5_) & (!g35) & (g14) & (g85)) + ((!i_3_) & (!i_5_) & (g35) & (!g14) & (!g85)) + ((!i_3_) & (!i_5_) & (g35) & (!g14) & (g85)) + ((!i_3_) & (!i_5_) & (g35) & (g14) & (!g85)) + ((!i_3_) & (!i_5_) & (g35) & (g14) & (g85)) + ((!i_3_) & (i_5_) & (!g35) & (g14) & (g85)) + ((!i_3_) & (i_5_) & (g35) & (g14) & (g85)) + ((i_3_) & (!i_5_) & (!g35) & (g14) & (g85)) + ((i_3_) & (!i_5_) & (g35) & (g14) & (g85)) + ((i_3_) & (i_5_) & (!g35) & (g14) & (g85)) + ((i_3_) & (i_5_) & (g35) & (g14) & (g85)));
	assign g298 = (((!g23) & (!g24) & (!g70) & (!g296) & (!g297)) + ((!g23) & (g24) & (!g70) & (!g296) & (!g297)) + ((!g23) & (g24) & (!g70) & (!g296) & (g297)) + ((g23) & (!g24) & (!g70) & (!g296) & (!g297)) + ((g23) & (!g24) & (g70) & (!g296) & (!g297)) + ((g23) & (g24) & (!g70) & (!g296) & (!g297)) + ((g23) & (g24) & (!g70) & (!g296) & (g297)) + ((g23) & (g24) & (g70) & (!g296) & (!g297)) + ((g23) & (g24) & (g70) & (!g296) & (g297)));
	assign g299 = (((!g292) & (!g293) & (g295) & (g298)));
	assign g302 = (((!i_6_) & (!g21) & (!g1) & (g137) & (!g59)) + ((!i_6_) & (g21) & (!g1) & (g137) & (!g59)) + ((i_6_) & (!g21) & (!g1) & (g137) & (!g59)) + ((i_6_) & (!g21) & (!g1) & (g137) & (g59)) + ((i_6_) & (g21) & (!g1) & (g137) & (!g59)));
	assign g303 = (((!g27) & (!g63) & (!g38) & (!g96)) + ((!g27) & (!g63) & (g38) & (!g96)) + ((!g27) & (g63) & (g38) & (!g96)) + ((g27) & (!g63) & (!g38) & (!g96)) + ((g27) & (!g63) & (g38) & (!g96)) + ((g27) & (g63) & (!g38) & (!g96)) + ((g27) & (g63) & (g38) & (!g96)));
	assign g304 = (((!g35) & (!g45) & (!g13) & (g4) & (!g243)) + ((!g35) & (!g45) & (!g13) & (g4) & (g243)) + ((!g35) & (g45) & (!g13) & (g4) & (!g243)) + ((!g35) & (g45) & (!g13) & (g4) & (g243)) + ((g35) & (!g45) & (!g13) & (!g4) & (!g243)) + ((g35) & (!g45) & (!g13) & (!g4) & (g243)) + ((g35) & (!g45) & (!g13) & (g4) & (!g243)) + ((g35) & (!g45) & (!g13) & (g4) & (g243)) + ((g35) & (!g45) & (g13) & (!g4) & (g243)) + ((g35) & (!g45) & (g13) & (g4) & (g243)) + ((g35) & (g45) & (!g13) & (!g4) & (g243)) + ((g35) & (g45) & (!g13) & (g4) & (!g243)) + ((g35) & (g45) & (!g13) & (g4) & (g243)) + ((g35) & (g45) & (g13) & (!g4) & (g243)) + ((g35) & (g45) & (g13) & (g4) & (g243)));
	assign g305 = (((!g2) & (g6) & (!g75) & (g71)) + ((!g2) & (g6) & (g75) & (g71)) + ((g2) & (!g6) & (g75) & (!g71)) + ((g2) & (!g6) & (g75) & (g71)) + ((g2) & (g6) & (!g75) & (g71)) + ((g2) & (g6) & (g75) & (!g71)) + ((g2) & (g6) & (g75) & (g71)));
	assign g306 = (((!g23) & (!g184) & (!g304) & (g607) & (!g305)) + ((g23) & (!g184) & (!g304) & (g607) & (!g305)) + ((g23) & (g184) & (!g304) & (g607) & (!g305)));
	assign g308 = (((!i_3_) & (!i_4_) & (!i_0_) & (i_2_) & (!g12) & (g219)) + ((!i_3_) & (!i_4_) & (!i_0_) & (i_2_) & (g12) & (g219)) + ((!i_3_) & (!i_4_) & (i_0_) & (i_2_) & (!g12) & (g219)) + ((!i_3_) & (!i_4_) & (i_0_) & (i_2_) & (g12) & (g219)) + ((!i_3_) & (i_4_) & (!i_0_) & (i_2_) & (!g12) & (g219)) + ((!i_3_) & (i_4_) & (!i_0_) & (i_2_) & (g12) & (g219)) + ((!i_3_) & (i_4_) & (i_0_) & (i_2_) & (!g12) & (g219)) + ((!i_3_) & (i_4_) & (i_0_) & (i_2_) & (g12) & (g219)) + ((i_3_) & (!i_4_) & (!i_0_) & (i_2_) & (g12) & (!g219)) + ((i_3_) & (!i_4_) & (!i_0_) & (i_2_) & (g12) & (g219)));
	assign g309 = (((!g42) & (!g23) & (!g194) & (g98)) + ((!g42) & (!g23) & (g194) & (g98)) + ((g42) & (!g23) & (!g194) & (g98)) + ((g42) & (!g23) & (g194) & (!g98)) + ((g42) & (!g23) & (g194) & (g98)) + ((g42) & (g23) & (g194) & (!g98)) + ((g42) & (g23) & (g194) & (g98)));
	assign g311 = (((!g2) & (!g23) & (!g59) & (!g13) & (g84)) + ((!g2) & (!g23) & (!g59) & (g13) & (g84)) + ((!g2) & (!g23) & (g59) & (!g13) & (g84)) + ((!g2) & (!g23) & (g59) & (g13) & (g84)) + ((g2) & (!g23) & (!g59) & (!g13) & (!g84)) + ((g2) & (!g23) & (!g59) & (!g13) & (g84)) + ((g2) & (!g23) & (!g59) & (g13) & (g84)) + ((g2) & (!g23) & (g59) & (!g13) & (g84)) + ((g2) & (!g23) & (g59) & (g13) & (g84)) + ((g2) & (g23) & (!g59) & (!g13) & (!g84)) + ((g2) & (g23) & (!g59) & (!g13) & (g84)));
	assign g316 = (((!g6) & (!g105) & (!g315)) + ((!g6) & (g105) & (!g315)) + ((g6) & (g105) & (!g315)));
	assign g317 = (((!g48) & (!g313) & (!g314) & (!g52) & (g316)) + ((!g48) & (!g313) & (!g314) & (g52) & (g316)) + ((g48) & (!g313) & (!g314) & (!g52) & (g316)));
	assign g318 = (((!g168) & (g310) & (g312) & (g317)));
	assign g319 = (((!g301) & (g211) & (g307) & (!g308) & (g318)));
	assign g320 = (((g90) & (g224) & (g274) & (g618) & (g300) & (g319)));
	assign g321 = (((!i_6_) & (i_7_) & (!i_8_) & (!g26) & (g243) & (!g268)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g26) & (g243) & (g268)) + ((!i_6_) & (i_7_) & (!i_8_) & (g26) & (g243) & (!g268)) + ((!i_6_) & (i_7_) & (!i_8_) & (g26) & (g243) & (g268)) + ((!i_6_) & (i_7_) & (i_8_) & (!g26) & (!g243) & (g268)) + ((!i_6_) & (i_7_) & (i_8_) & (!g26) & (g243) & (g268)) + ((!i_6_) & (i_7_) & (i_8_) & (g26) & (!g243) & (g268)) + ((!i_6_) & (i_7_) & (i_8_) & (g26) & (g243) & (g268)) + ((i_6_) & (!i_7_) & (!i_8_) & (g26) & (!g243) & (!g268)) + ((i_6_) & (!i_7_) & (!i_8_) & (g26) & (!g243) & (g268)) + ((i_6_) & (!i_7_) & (!i_8_) & (g26) & (g243) & (!g268)) + ((i_6_) & (!i_7_) & (!i_8_) & (g26) & (g243) & (g268)) + ((i_6_) & (i_7_) & (!i_8_) & (!g26) & (g243) & (!g268)) + ((i_6_) & (i_7_) & (!i_8_) & (!g26) & (g243) & (g268)) + ((i_6_) & (i_7_) & (!i_8_) & (g26) & (g243) & (!g268)) + ((i_6_) & (i_7_) & (!i_8_) & (g26) & (g243) & (g268)) + ((i_6_) & (i_7_) & (i_8_) & (!g26) & (!g243) & (g268)) + ((i_6_) & (i_7_) & (i_8_) & (!g26) & (g243) & (g268)) + ((i_6_) & (i_7_) & (i_8_) & (g26) & (!g243) & (g268)) + ((i_6_) & (i_7_) & (i_8_) & (g26) & (g243) & (g268)));
	assign g322 = (((!g27) & (!g45) & (!g1) & (!g6) & (g16)) + ((!g27) & (!g45) & (!g1) & (g6) & (!g16)) + ((!g27) & (!g45) & (!g1) & (g6) & (g16)) + ((!g27) & (!g45) & (g1) & (g6) & (!g16)) + ((!g27) & (!g45) & (g1) & (g6) & (g16)) + ((!g27) & (g45) & (!g1) & (!g6) & (g16)) + ((!g27) & (g45) & (!g1) & (g6) & (g16)) + ((g27) & (!g45) & (!g1) & (!g6) & (g16)) + ((g27) & (!g45) & (!g1) & (g6) & (g16)) + ((g27) & (g45) & (!g1) & (!g6) & (g16)) + ((g27) & (g45) & (!g1) & (g6) & (g16)));
	assign g324 = (((!g28) & (g48) & (!g189) & (g184)) + ((!g28) & (g48) & (g189) & (g184)) + ((g28) & (!g48) & (g189) & (!g184)) + ((g28) & (!g48) & (g189) & (g184)) + ((g28) & (g48) & (!g189) & (g184)) + ((g28) & (g48) & (g189) & (!g184)) + ((g28) & (g48) & (g189) & (g184)));
	assign g325 = (((g137) & (g134) & (g230)));
	assign g326 = (((!g35) & (!g25) & (!g59) & (!g4) & (!g325)) + ((!g35) & (!g25) & (g59) & (!g4) & (!g325)) + ((!g35) & (g25) & (!g59) & (!g4) & (!g325)) + ((!g35) & (g25) & (!g59) & (g4) & (!g325)) + ((!g35) & (g25) & (g59) & (!g4) & (!g325)) + ((!g35) & (g25) & (g59) & (g4) & (!g325)) + ((g35) & (!g25) & (g59) & (!g4) & (!g325)) + ((g35) & (g25) & (!g59) & (!g4) & (!g325)) + ((g35) & (g25) & (!g59) & (g4) & (!g325)) + ((g35) & (g25) & (g59) & (!g4) & (!g325)) + ((g35) & (g25) & (g59) & (g4) & (!g325)));
	assign g328 = (((!i_6_) & (g14) & (g26) & (!g99)) + ((!i_6_) & (g14) & (g26) & (g99)) + ((i_6_) & (g14) & (!g26) & (g99)) + ((i_6_) & (g14) & (g26) & (g99)));
	assign g329 = (((!g45) & (!g6) & (!g24) & (g67) & (!g91)) + ((!g45) & (!g6) & (!g24) & (g67) & (g91)) + ((!g45) & (!g6) & (g24) & (g67) & (!g91)) + ((!g45) & (!g6) & (g24) & (g67) & (g91)) + ((!g45) & (g6) & (!g24) & (!g67) & (!g91)) + ((!g45) & (g6) & (!g24) & (!g67) & (g91)) + ((!g45) & (g6) & (!g24) & (g67) & (!g91)) + ((!g45) & (g6) & (!g24) & (g67) & (g91)) + ((!g45) & (g6) & (g24) & (!g67) & (g91)) + ((!g45) & (g6) & (g24) & (g67) & (!g91)) + ((!g45) & (g6) & (g24) & (g67) & (g91)) + ((g45) & (g6) & (!g24) & (!g67) & (g91)) + ((g45) & (g6) & (!g24) & (g67) & (g91)) + ((g45) & (g6) & (g24) & (!g67) & (g91)) + ((g45) & (g6) & (g24) & (g67) & (g91)));
	assign g331 = (((g14) & (g64) & (g230)));
	assign g333 = (((i_3_) & (!i_4_) & (!i_5_) & (!i_6_) & (i_7_) & (i_8_)) + ((i_3_) & (i_4_) & (i_5_) & (!i_6_) & (!i_7_) & (!i_8_)));
	assign g335 = (((!g11) & (!g35) & (!g28) & (!g25) & (!g38) & (!g334)) + ((!g11) & (!g35) & (!g28) & (!g25) & (g38) & (!g334)) + ((!g11) & (!g35) & (!g28) & (g25) & (!g38) & (!g334)) + ((!g11) & (!g35) & (!g28) & (g25) & (g38) & (!g334)) + ((!g11) & (!g35) & (g28) & (!g25) & (g38) & (!g334)) + ((!g11) & (!g35) & (g28) & (g25) & (!g38) & (!g334)) + ((!g11) & (!g35) & (g28) & (g25) & (g38) & (!g334)) + ((!g11) & (g35) & (!g28) & (g25) & (!g38) & (!g334)) + ((!g11) & (g35) & (!g28) & (g25) & (g38) & (!g334)) + ((!g11) & (g35) & (g28) & (g25) & (!g38) & (!g334)) + ((!g11) & (g35) & (g28) & (g25) & (g38) & (!g334)) + ((g11) & (!g35) & (!g28) & (!g25) & (!g38) & (!g334)) + ((g11) & (!g35) & (!g28) & (!g25) & (g38) & (!g334)) + ((g11) & (!g35) & (!g28) & (g25) & (!g38) & (!g334)) + ((g11) & (!g35) & (!g28) & (g25) & (g38) & (!g334)) + ((g11) & (!g35) & (g28) & (!g25) & (g38) & (!g334)) + ((g11) & (!g35) & (g28) & (g25) & (!g38) & (!g334)) + ((g11) & (!g35) & (g28) & (g25) & (g38) & (!g334)) + ((g11) & (g35) & (!g28) & (!g25) & (!g38) & (!g334)) + ((g11) & (g35) & (!g28) & (!g25) & (g38) & (!g334)) + ((g11) & (g35) & (!g28) & (g25) & (!g38) & (!g334)) + ((g11) & (g35) & (!g28) & (g25) & (g38) & (!g334)) + ((g11) & (g35) & (g28) & (!g25) & (g38) & (!g334)) + ((g11) & (g35) & (g28) & (g25) & (!g38) & (!g334)) + ((g11) & (g35) & (g28) & (g25) & (g38) & (!g334)));
	assign g336 = (((!i_3_) & (!g21) & (!g42) & (!g8) & (g7)) + ((!i_3_) & (!g21) & (!g42) & (g8) & (g7)) + ((!i_3_) & (!g21) & (g42) & (!g8) & (g7)) + ((!i_3_) & (!g21) & (g42) & (g8) & (g7)) + ((i_3_) & (!g21) & (!g42) & (!g8) & (g7)) + ((i_3_) & (!g21) & (!g42) & (g8) & (g7)) + ((i_3_) & (!g21) & (g42) & (!g8) & (g7)) + ((i_3_) & (!g21) & (g42) & (g8) & (!g7)) + ((i_3_) & (!g21) & (g42) & (g8) & (g7)) + ((i_3_) & (g21) & (g42) & (g8) & (!g7)) + ((i_3_) & (g21) & (g42) & (g8) & (g7)));
	assign g337 = (((!i_6_) & (i_7_) & (!i_8_) & (!g70) & (g184)) + ((!i_6_) & (i_7_) & (!i_8_) & (g70) & (g184)) + ((i_6_) & (!i_7_) & (!i_8_) & (g70) & (!g184)) + ((i_6_) & (!i_7_) & (!i_8_) & (g70) & (g184)) + ((i_6_) & (i_7_) & (!i_8_) & (!g70) & (g184)) + ((i_6_) & (i_7_) & (!i_8_) & (g70) & (g184)));
	assign g338 = (((g46) & (!g48) & (g60)) + ((g46) & (g48) & (!g60)) + ((g46) & (g48) & (g60)));
	assign g339 = (((!g2) & (!g98) & (!g252) & (!g337) & (!g338)) + ((!g2) & (g98) & (!g252) & (!g337) & (!g338)) + ((g2) & (!g98) & (!g252) & (!g337) & (!g338)));
	assign g340 = (((g312) & (g332) & (g335) & (!g336) & (g339)));
	assign g342 = (((!i_0_) & (!g27) & (g14) & (!g135) & (g217)) + ((!i_0_) & (!g27) & (g14) & (g135) & (g217)) + ((i_0_) & (!g27) & (!g14) & (g135) & (!g217)) + ((i_0_) & (!g27) & (!g14) & (g135) & (g217)) + ((i_0_) & (!g27) & (g14) & (!g135) & (g217)) + ((i_0_) & (!g27) & (g14) & (g135) & (!g217)) + ((i_0_) & (!g27) & (g14) & (g135) & (g217)) + ((i_0_) & (g27) & (!g14) & (g135) & (!g217)) + ((i_0_) & (g27) & (!g14) & (g135) & (g217)) + ((i_0_) & (g27) & (g14) & (g135) & (!g217)) + ((i_0_) & (g27) & (g14) & (g135) & (g217)));
	assign g345 = (((!i_5_) & (i_6_) & (!i_7_) & (!i_8_) & (g5)) + ((!i_5_) & (i_6_) & (i_7_) & (!i_8_) & (g5)) + ((i_5_) & (!i_6_) & (i_7_) & (!i_8_) & (g5)));
	assign g347 = (((!i_6_) & (!i_7_) & (!i_8_) & (g46) & (!g77) & (!g189)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g46) & (!g77) & (g189)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g46) & (g77) & (!g189)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g46) & (g77) & (g189)) + ((i_6_) & (!i_7_) & (!i_8_) & (g46) & (!g77) & (!g189)) + ((i_6_) & (!i_7_) & (!i_8_) & (g46) & (!g77) & (g189)) + ((i_6_) & (!i_7_) & (!i_8_) & (g46) & (g77) & (!g189)) + ((i_6_) & (!i_7_) & (!i_8_) & (g46) & (g77) & (g189)) + ((i_6_) & (!i_7_) & (i_8_) & (!g46) & (!g77) & (g189)) + ((i_6_) & (!i_7_) & (i_8_) & (!g46) & (g77) & (!g189)) + ((i_6_) & (!i_7_) & (i_8_) & (!g46) & (g77) & (g189)) + ((i_6_) & (!i_7_) & (i_8_) & (g46) & (!g77) & (g189)) + ((i_6_) & (!i_7_) & (i_8_) & (g46) & (g77) & (!g189)) + ((i_6_) & (!i_7_) & (i_8_) & (g46) & (g77) & (g189)) + ((i_6_) & (i_7_) & (!i_8_) & (g46) & (!g77) & (!g189)) + ((i_6_) & (i_7_) & (!i_8_) & (g46) & (!g77) & (g189)) + ((i_6_) & (i_7_) & (!i_8_) & (g46) & (g77) & (!g189)) + ((i_6_) & (i_7_) & (!i_8_) & (g46) & (g77) & (g189)));
	assign g348 = (((i_3_) & (!i_4_) & (i_0_) & (!i_1_)));
	assign g349 = (((!g2) & (!g161) & (!g296) & (!g348)) + ((!g2) & (!g161) & (!g296) & (g348)) + ((!g2) & (g161) & (!g296) & (!g348)) + ((!g2) & (g161) & (!g296) & (g348)) + ((g2) & (!g161) & (!g296) & (!g348)));
	assign g350 = (((g343) & (!g344) & (!g346) & (!g347) & (g349)));
	assign g351 = (((!i_5_) & (!i_2_) & (!g48) & (!g219)) + ((!i_5_) & (i_2_) & (!g48) & (!g219)) + ((!i_5_) & (i_2_) & (g48) & (!g219)) + ((i_5_) & (!i_2_) & (!g48) & (!g219)) + ((i_5_) & (!i_2_) & (g48) & (!g219)) + ((i_5_) & (i_2_) & (!g48) & (!g219)) + ((i_5_) & (i_2_) & (g48) & (!g219)));
	assign g353 = (((g50) & (i_6_) & (!i_7_) & (g86)));
	assign g354 = (((!g13) & (!g4) & (!g352) & (g125) & (!g353)) + ((g13) & (!g4) & (!g352) & (g125) & (!g353)) + ((g13) & (g4) & (!g352) & (g125) & (!g353)));
	assign g355 = (((!g301) & (g20) & (!g342) & (g350) & (g354)));
	assign g356 = (((g178) & (g234) & (g323) & (g341) & (g355)));
	assign g357 = (((!g6) & (g4) & (g110) & (!g243)) + ((!g6) & (g4) & (g110) & (g243)) + ((g6) & (!g4) & (!g110) & (g243)) + ((g6) & (!g4) & (g110) & (g243)) + ((g6) & (g4) & (!g110) & (g243)) + ((g6) & (g4) & (g110) & (!g243)) + ((g6) & (g4) & (g110) & (g243)));
	assign g360 = (((!i_6_) & (!i_7_) & (!i_8_) & (!g73) & (!g184) & (g359)) + ((!i_6_) & (!i_7_) & (!i_8_) & (!g73) & (g184) & (g359)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g73) & (!g184) & (g359)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g73) & (g184) & (g359)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g73) & (g184) & (!g359)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g73) & (g184) & (g359)) + ((!i_6_) & (!i_7_) & (i_8_) & (g73) & (!g184) & (!g359)) + ((!i_6_) & (!i_7_) & (i_8_) & (g73) & (!g184) & (g359)) + ((!i_6_) & (!i_7_) & (i_8_) & (g73) & (g184) & (!g359)) + ((!i_6_) & (!i_7_) & (i_8_) & (g73) & (g184) & (g359)) + ((i_6_) & (!i_7_) & (i_8_) & (g73) & (!g184) & (!g359)) + ((i_6_) & (!i_7_) & (i_8_) & (g73) & (!g184) & (g359)) + ((i_6_) & (!i_7_) & (i_8_) & (g73) & (g184) & (!g359)) + ((i_6_) & (!i_7_) & (i_8_) & (g73) & (g184) & (g359)));
	assign g361 = (((g127) & (!i_2_) & (!i_6_) & (g137) & (g5)) + ((g127) & (i_2_) & (i_6_) & (g137) & (g5)));
	assign g362 = (((!g11) & (!g42) & (!g22) & (!g121) & (!g361)) + ((!g11) & (!g42) & (g22) & (!g121) & (!g361)) + ((!g11) & (g42) & (!g22) & (!g121) & (!g361)) + ((g11) & (!g42) & (!g22) & (!g121) & (!g361)) + ((g11) & (!g42) & (!g22) & (g121) & (!g361)) + ((g11) & (!g42) & (g22) & (!g121) & (!g361)) + ((g11) & (!g42) & (g22) & (g121) & (!g361)) + ((g11) & (g42) & (!g22) & (!g121) & (!g361)) + ((g11) & (g42) & (!g22) & (g121) & (!g361)));
	assign g365 = (((!g21) & (!g38) & (!g7) & (!g265) & (!g364)) + ((!g21) & (g38) & (!g7) & (!g265) & (!g364)) + ((!g21) & (g38) & (g7) & (!g265) & (!g364)) + ((g21) & (!g38) & (!g7) & (!g265) & (!g364)) + ((g21) & (!g38) & (!g7) & (g265) & (!g364)) + ((g21) & (g38) & (!g7) & (!g265) & (!g364)) + ((g21) & (g38) & (!g7) & (g265) & (!g364)) + ((g21) & (g38) & (g7) & (!g265) & (!g364)) + ((g21) & (g38) & (g7) & (g265) & (!g364)));
	assign g366 = (((!g175) & (!g256) & (!g363) & (g365)));
	assign g369 = (((!g50) & (i_6_) & (g14) & (!g25) & (g129)) + ((!g50) & (i_6_) & (g14) & (g25) & (g129)) + ((g50) & (i_6_) & (g14) & (!g25) & (!g129)) + ((g50) & (i_6_) & (g14) & (!g25) & (g129)) + ((g50) & (i_6_) & (g14) & (g25) & (g129)));
	assign g370 = (((!i_6_) & (!g45) & (!g1) & (g47) & (!g110)) + ((!i_6_) & (!g45) & (!g1) & (g47) & (g110)) + ((i_6_) & (!g45) & (!g1) & (g47) & (g110)) + ((i_6_) & (!g45) & (g1) & (g47) & (g110)));
	assign g372 = (((!i_6_) & (!i_7_) & (!i_8_) & (g77) & (!g99)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g77) & (g99)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g77) & (g99)) + ((!i_6_) & (!i_7_) & (i_8_) & (g77) & (g99)) + ((i_6_) & (!i_7_) & (i_8_) & (g77) & (!g99)) + ((i_6_) & (!i_7_) & (i_8_) & (g77) & (g99)));
	assign g373 = (((!g67) & (!g116) & (!g290)) + ((!g67) & (g116) & (!g290)) + ((g67) & (!g116) & (!g290)));
	assign g374 = (((!g173) & (!g294) & (!g145) & (g140) & (g373)));
	assign g375 = (((!g23) & (!g75) & (!g160) & (!g372) & (g374)) + ((g23) & (!g75) & (!g160) & (!g372) & (g374)) + ((g23) & (g75) & (!g160) & (!g372) & (g374)));
	assign g377 = (((!i_6_) & (!i_7_) & (!i_8_) & (!g24) & (!g64) & (g26)) + ((!i_6_) & (!i_7_) & (!i_8_) & (!g24) & (g64) & (g26)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g24) & (!g64) & (g26)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g24) & (g64) & (g26)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g24) & (!g64) & (g26)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g24) & (g64) & (g26)) + ((!i_6_) & (i_7_) & (!i_8_) & (g24) & (!g64) & (g26)) + ((!i_6_) & (i_7_) & (!i_8_) & (g24) & (g64) & (g26)) + ((!i_6_) & (i_7_) & (i_8_) & (!g24) & (g64) & (!g26)) + ((!i_6_) & (i_7_) & (i_8_) & (!g24) & (g64) & (g26)) + ((i_6_) & (i_7_) & (i_8_) & (!g24) & (g64) & (!g26)) + ((i_6_) & (i_7_) & (i_8_) & (!g24) & (g64) & (g26)));
	assign g378 = (((!g204) & (!g376) & (g246) & (g249) & (!g377)));
	assign g379 = (((!i_0_) & (!i_1_) & (i_2_) & (!g23) & (g123)) + ((!i_0_) & (!i_1_) & (i_2_) & (g23) & (g123)) + ((!i_0_) & (i_1_) & (i_2_) & (!g23) & (g123)) + ((!i_0_) & (i_1_) & (i_2_) & (g23) & (g123)) + ((i_0_) & (!i_1_) & (i_2_) & (!g23) & (!g123)) + ((i_0_) & (!i_1_) & (i_2_) & (!g23) & (g123)));
	assign g380 = (((!i_3_) & (!g195) & (!g379) & (g90) & (g618)) + ((i_3_) & (!g195) & (!g379) & (g90) & (g618)) + ((i_3_) & (!g195) & (g379) & (g90) & (g618)));
	assign g382 = (((!i_6_) & (g63) & (!g21) & (!g25) & (!g110) & (!g218)) + ((!i_6_) & (g63) & (!g21) & (!g25) & (!g110) & (g218)) + ((!i_6_) & (g63) & (!g21) & (!g25) & (g110) & (!g218)) + ((!i_6_) & (g63) & (!g21) & (!g25) & (g110) & (g218)) + ((!i_6_) & (g63) & (!g21) & (g25) & (!g110) & (g218)) + ((!i_6_) & (g63) & (!g21) & (g25) & (g110) & (g218)) + ((!i_6_) & (g63) & (g21) & (!g25) & (!g110) & (g218)) + ((!i_6_) & (g63) & (g21) & (!g25) & (g110) & (g218)) + ((!i_6_) & (g63) & (g21) & (g25) & (!g110) & (g218)) + ((!i_6_) & (g63) & (g21) & (g25) & (g110) & (g218)) + ((i_6_) & (g63) & (!g21) & (!g25) & (!g110) & (g218)) + ((i_6_) & (g63) & (!g21) & (!g25) & (g110) & (!g218)) + ((i_6_) & (g63) & (!g21) & (!g25) & (g110) & (g218)) + ((i_6_) & (g63) & (!g21) & (g25) & (!g110) & (g218)) + ((i_6_) & (g63) & (!g21) & (g25) & (g110) & (!g218)) + ((i_6_) & (g63) & (!g21) & (g25) & (g110) & (g218)) + ((i_6_) & (g63) & (g21) & (!g25) & (!g110) & (g218)) + ((i_6_) & (g63) & (g21) & (!g25) & (g110) & (g218)) + ((i_6_) & (g63) & (g21) & (g25) & (!g110) & (g218)) + ((i_6_) & (g63) & (g21) & (g25) & (g110) & (g218)));
	assign g385 = (((!g27) & (!g21) & (!g6) & (!g3) & (g121)) + ((!g27) & (!g21) & (!g6) & (g3) & (g121)) + ((!g27) & (!g21) & (g6) & (!g3) & (g121)) + ((!g27) & (!g21) & (g6) & (g3) & (!g121)) + ((!g27) & (!g21) & (g6) & (g3) & (g121)) + ((!g27) & (g21) & (g6) & (g3) & (!g121)) + ((!g27) & (g21) & (g6) & (g3) & (g121)) + ((g27) & (!g21) & (!g6) & (!g3) & (g121)) + ((g27) & (!g21) & (!g6) & (g3) & (g121)) + ((g27) & (!g21) & (g6) & (!g3) & (g121)) + ((g27) & (!g21) & (g6) & (g3) & (g121)));
	assign g388 = (((!g1) & (!g159) & (!g150) & (!g387)) + ((g1) & (!g159) & (!g150) & (!g387)) + ((g1) & (g159) & (!g150) & (!g387)));
	assign g390 = (((!g18) & (!g170) & (!g389)));
	assign g391 = (((g127) & (!i_2_) & (!i_6_) & (i_7_) & (!i_8_) & (g3)) + ((g127) & (!i_2_) & (i_6_) & (!i_7_) & (!i_8_) & (g3)) + ((g127) & (!i_2_) & (i_6_) & (!i_7_) & (i_8_) & (g3)) + ((g127) & (!i_2_) & (i_6_) & (i_7_) & (!i_8_) & (g3)) + ((g127) & (i_2_) & (!i_6_) & (i_7_) & (!i_8_) & (g3)) + ((g127) & (i_2_) & (i_6_) & (i_7_) & (!i_8_) & (g3)));
	assign g393 = (((!g344) & (g388) & (g390) & (!g391) & (g583)));
	assign g394 = (((!g72) & (g166) & (g383) & (g386) & (g393)));
	assign g395 = (((g274) & (g283) & (g367) & (g381) & (g394)));
	assign g397 = (((!i_4_) & (!g42) & (!g12) & (g9)) + ((!i_4_) & (!g42) & (g12) & (g9)) + ((!i_4_) & (g42) & (!g12) & (g9)) + ((!i_4_) & (g42) & (g12) & (g9)) + ((i_4_) & (g42) & (g12) & (!g9)) + ((i_4_) & (g42) & (g12) & (g9)));
	assign g399 = (((!g21) & (!g42) & (!g12) & (!g75) & (!g124)) + ((!g21) & (!g42) & (!g12) & (g75) & (!g124)) + ((!g21) & (!g42) & (g12) & (!g75) & (!g124)) + ((!g21) & (g42) & (!g12) & (!g75) & (!g124)) + ((!g21) & (g42) & (!g12) & (g75) & (!g124)) + ((g21) & (!g42) & (!g12) & (!g75) & (!g124)) + ((g21) & (!g42) & (!g12) & (g75) & (!g124)) + ((g21) & (!g42) & (g12) & (!g75) & (!g124)) + ((g21) & (g42) & (!g12) & (!g75) & (!g124)) + ((g21) & (g42) & (!g12) & (g75) & (!g124)) + ((g21) & (g42) & (g12) & (!g75) & (!g124)));
	assign g403 = (((!i_6_) & (!i_7_) & (i_8_) & (!g77) & (g71) & (!g161)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g77) & (g71) & (g161)) + ((!i_6_) & (!i_7_) & (i_8_) & (g77) & (g71) & (!g161)) + ((!i_6_) & (!i_7_) & (i_8_) & (g77) & (g71) & (g161)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g77) & (!g71) & (g161)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g77) & (g71) & (!g161)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g77) & (g71) & (g161)) + ((i_6_) & (!i_7_) & (!i_8_) & (g77) & (!g71) & (g161)) + ((i_6_) & (!i_7_) & (!i_8_) & (g77) & (g71) & (!g161)) + ((i_6_) & (!i_7_) & (!i_8_) & (g77) & (g71) & (g161)) + ((i_6_) & (i_7_) & (i_8_) & (g77) & (!g71) & (!g161)) + ((i_6_) & (i_7_) & (i_8_) & (g77) & (!g71) & (g161)) + ((i_6_) & (i_7_) & (i_8_) & (g77) & (g71) & (!g161)) + ((i_6_) & (i_7_) & (i_8_) & (g77) & (g71) & (g161)));
	assign g404 = (((!g402) & (g93) & (g631) & (!g403)));
	assign g407 = (((!g50) & (g48) & (g88) & (!g111) & (!g230)) + ((!g50) & (g48) & (g88) & (!g111) & (g230)) + ((!g50) & (g48) & (g88) & (g111) & (!g230)) + ((!g50) & (g48) & (g88) & (g111) & (g230)) + ((g50) & (!g48) & (!g88) & (g111) & (g230)) + ((g50) & (!g48) & (g88) & (g111) & (g230)) + ((g50) & (g48) & (!g88) & (g111) & (g230)) + ((g50) & (g48) & (g88) & (!g111) & (!g230)) + ((g50) & (g48) & (g88) & (!g111) & (g230)) + ((g50) & (g48) & (g88) & (g111) & (!g230)) + ((g50) & (g48) & (g88) & (g111) & (g230)));
	assign g410 = (((!g35) & (!g48) & (!g117) & (!g334)) + ((!g35) & (!g48) & (g117) & (!g334)) + ((!g35) & (g48) & (!g117) & (!g334)) + ((g35) & (!g48) & (!g117) & (!g334)) + ((g35) & (g48) & (!g117) & (!g334)));
	assign g411 = (((!i_4_) & (!i_5_) & (!i_0_) & (i_1_) & (g12)));
	assign g412 = (((!g8) & (!g137) & (!g91) & (!g243) & (!g411)) + ((!g8) & (!g137) & (!g91) & (g243) & (!g411)) + ((!g8) & (!g137) & (g91) & (!g243) & (!g411)) + ((!g8) & (!g137) & (g91) & (g243) & (!g411)) + ((!g8) & (g137) & (!g91) & (!g243) & (!g411)) + ((!g8) & (g137) & (g91) & (!g243) & (!g411)) + ((g8) & (!g137) & (!g91) & (!g243) & (!g411)) + ((g8) & (!g137) & (!g91) & (g243) & (!g411)) + ((g8) & (g137) & (!g91) & (!g243) & (!g411)));
	assign g414 = (((!i_5_) & (!g6) & (g5) & (g110) & (g111)) + ((!i_5_) & (g6) & (g5) & (g110) & (!g111)) + ((!i_5_) & (g6) & (g5) & (g110) & (g111)) + ((i_5_) & (g6) & (g5) & (g110) & (!g111)) + ((i_5_) & (g6) & (g5) & (g110) & (g111)));
	assign g415 = (((!g23) & (!g359) & (!g413) & (!g414)) + ((g23) & (!g359) & (!g413) & (!g414)) + ((g23) & (g359) & (!g413) & (!g414)));
	assign g416 = (((!g87) & (!g346) & (g410) & (g412) & (g415)));
	assign g417 = (((g254) & (g307) & (g289) & (!g409) & (g416)));
	assign g418 = (((g381) & (g405) & (g408) & (g417)));
	assign g420 = (((!i_0_) & (!i_1_) & (i_2_) & (!i_6_) & (i_7_) & (i_8_)) + ((!i_0_) & (i_1_) & (!i_2_) & (!i_6_) & (!i_7_) & (!i_8_)) + ((!i_0_) & (i_1_) & (!i_2_) & (!i_6_) & (!i_7_) & (i_8_)));
	assign g421 = (((!i_0_) & (!i_6_) & (!g38) & (g420)));
	assign g422 = (((g28) & (!g42) & (!g45) & (!g1) & (g32)) + ((g28) & (!g42) & (g45) & (!g1) & (g32)) + ((g28) & (g42) & (!g45) & (!g1) & (!g32)) + ((g28) & (g42) & (!g45) & (!g1) & (g32)) + ((g28) & (g42) & (!g45) & (g1) & (!g32)) + ((g28) & (g42) & (!g45) & (g1) & (g32)) + ((g28) & (g42) & (g45) & (!g1) & (g32)));
	assign g423 = (((!g27) & (!g6) & (!g36) & (!g422) & (g572)) + ((!g27) & (!g6) & (g36) & (!g422) & (g572)) + ((!g27) & (g6) & (g36) & (!g422) & (g572)) + ((g27) & (!g6) & (!g36) & (!g422) & (g572)) + ((g27) & (!g6) & (g36) & (!g422) & (g572)) + ((g27) & (g6) & (!g36) & (!g422) & (g572)) + ((g27) & (g6) & (g36) & (!g422) & (g572)));
	assign g425 = (((!i_6_) & (!i_8_) & (!g21) & (!g1)));
	assign g426 = (((!i_6_) & (g14) & (g32) & (g110)) + ((i_6_) & (!g14) & (g32) & (g110)) + ((i_6_) & (g14) & (g32) & (g110)));
	assign g429 = (((!g11) & (!g29) & (!g428)) + ((g11) & (!g29) & (!g428)) + ((g11) & (g29) & (!g428)));
	assign g430 = (((!g63) & (!g45) & (!g129) & (g141)) + ((!g63) & (!g45) & (g129) & (g141)) + ((g63) & (!g45) & (!g129) & (g141)) + ((g63) & (!g45) & (g129) & (!g141)) + ((g63) & (!g45) & (g129) & (g141)) + ((g63) & (g45) & (g129) & (!g141)) + ((g63) & (g45) & (g129) & (g141)));
	assign g432 = (((!i_7_) & (!g8) & (!g25) & (!g32) & (!g97) & (!g217)) + ((!i_7_) & (!g8) & (!g25) & (!g32) & (!g97) & (g217)) + ((!i_7_) & (!g8) & (!g25) & (g32) & (!g97) & (!g217)) + ((!i_7_) & (!g8) & (!g25) & (g32) & (!g97) & (g217)) + ((!i_7_) & (!g8) & (g25) & (!g32) & (!g97) & (!g217)) + ((!i_7_) & (!g8) & (g25) & (!g32) & (!g97) & (g217)) + ((!i_7_) & (!g8) & (g25) & (g32) & (!g97) & (!g217)) + ((!i_7_) & (!g8) & (g25) & (g32) & (!g97) & (g217)) + ((!i_7_) & (g8) & (!g25) & (!g32) & (!g97) & (!g217)) + ((!i_7_) & (g8) & (!g25) & (!g32) & (!g97) & (g217)) + ((!i_7_) & (g8) & (g25) & (!g32) & (!g97) & (!g217)) + ((!i_7_) & (g8) & (g25) & (!g32) & (!g97) & (g217)) + ((!i_7_) & (g8) & (g25) & (g32) & (!g97) & (!g217)) + ((!i_7_) & (g8) & (g25) & (g32) & (!g97) & (g217)) + ((i_7_) & (!g8) & (!g25) & (!g32) & (!g97) & (!g217)) + ((i_7_) & (!g8) & (!g25) & (g32) & (!g97) & (!g217)) + ((i_7_) & (!g8) & (g25) & (!g32) & (!g97) & (!g217)) + ((i_7_) & (!g8) & (g25) & (!g32) & (!g97) & (g217)) + ((i_7_) & (!g8) & (g25) & (g32) & (!g97) & (!g217)) + ((i_7_) & (!g8) & (g25) & (g32) & (!g97) & (g217)) + ((i_7_) & (g8) & (!g25) & (!g32) & (!g97) & (!g217)) + ((i_7_) & (g8) & (g25) & (!g32) & (!g97) & (!g217)) + ((i_7_) & (g8) & (g25) & (!g32) & (!g97) & (g217)) + ((i_7_) & (g8) & (g25) & (g32) & (!g97) & (!g217)) + ((i_7_) & (g8) & (g25) & (g32) & (!g97) & (g217)));
	assign g433 = (((!i_1_) & (g6) & (g33) & (!g38)) + ((!i_1_) & (g6) & (g33) & (g38)) + ((i_1_) & (g6) & (!g33) & (!g38)) + ((i_1_) & (g6) & (g33) & (!g38)) + ((i_1_) & (g6) & (g33) & (g38)));
	assign g434 = (((!g35) & (!g189) & (!g229) & (!g431) & (g432) & (!g433)) + ((!g35) & (g189) & (!g229) & (!g431) & (g432) & (!g433)) + ((g35) & (!g189) & (!g229) & (!g431) & (g432) & (!g433)));
	assign g435 = (((!g352) & (g332) & (g429) & (!g430) & (g434)));
	assign g436 = (((!g419) & (g367) & (g424) & (g427) & (g435)));
	assign g437 = (((g31) & (g300) & (g371) & (g405) & (g436)));
	assign g439 = (((!g21) & (!g1) & (g2) & (!g24) & (!g36)) + ((!g21) & (!g1) & (g2) & (!g24) & (g36)) + ((!g21) & (!g1) & (g2) & (g24) & (!g36)) + ((!g21) & (g1) & (g2) & (!g24) & (!g36)) + ((!g21) & (g1) & (g2) & (!g24) & (g36)) + ((g21) & (!g1) & (g2) & (!g24) & (!g36)) + ((g21) & (!g1) & (g2) & (g24) & (!g36)));
	assign g441 = (((g137) & (g15) & (g440)));
	assign g442 = (((!g6) & (!g5) & (!g110) & (!g99) & (!g441)) + ((!g6) & (!g5) & (!g110) & (g99) & (!g441)) + ((!g6) & (!g5) & (g110) & (!g99) & (!g441)) + ((!g6) & (!g5) & (g110) & (g99) & (!g441)) + ((!g6) & (g5) & (!g110) & (!g99) & (!g441)) + ((!g6) & (g5) & (!g110) & (g99) & (!g441)) + ((!g6) & (g5) & (g110) & (!g99) & (!g441)) + ((!g6) & (g5) & (g110) & (g99) & (!g441)) + ((g6) & (!g5) & (!g110) & (!g99) & (!g441)) + ((g6) & (!g5) & (g110) & (!g99) & (!g441)) + ((g6) & (g5) & (!g110) & (!g99) & (!g441)));
	assign g443 = (((!g35) & (!g161) & (!g376) & (!g439) & (g442)) + ((!g35) & (g161) & (!g376) & (!g439) & (g442)) + ((g35) & (!g161) & (!g376) & (!g439) & (g442)));
	assign g444 = (((!i_8_) & (!g65) & (!g247) & (g398)) + ((!i_8_) & (g65) & (!g247) & (g398)) + ((i_8_) & (!g65) & (!g247) & (g398)));
	assign g446 = (((i_3_) & (i_1_) & (!i_2_) & (i_7_) & (g64)));
	assign g450 = (((!g255) & (!g384) & (g310) & (g559)));
	assign g451 = (((!g50) & (i_6_) & (i_8_) & (g5) & (!g13) & (!g17)) + ((!g50) & (i_6_) & (i_8_) & (g5) & (!g13) & (g17)) + ((g50) & (!i_6_) & (i_8_) & (!g5) & (!g13) & (g17)) + ((g50) & (!i_6_) & (i_8_) & (!g5) & (g13) & (g17)) + ((g50) & (!i_6_) & (i_8_) & (g5) & (!g13) & (g17)) + ((g50) & (!i_6_) & (i_8_) & (g5) & (g13) & (g17)) + ((g50) & (i_6_) & (i_8_) & (g5) & (!g13) & (!g17)) + ((g50) & (i_6_) & (i_8_) & (g5) & (!g13) & (g17)));
	assign g452 = (((!g275) & (!g402) & (g670) & (g147) & (!g451)));
	assign g453 = (((g80) & (g291) & (g383) & (g427) & (g450) & (g452)));
	assign g454 = (((g109) & (g341) & (g408) & (g445) & (g453)));
	assign g455 = (((g127) & (!i_2_) & (g2) & (!g60) & (!g38)) + ((g127) & (!i_2_) & (g2) & (g60) & (!g38)) + ((g127) & (i_2_) & (!g2) & (g60) & (!g38)) + ((g127) & (i_2_) & (g2) & (g60) & (!g38)));
	assign g459 = (((!g267) & (!g313) & (!g389) & (!g419) & (!g457) & (!g458)));
	assign g460 = (((!i_4_) & (i_5_) & (i_1_) & (i_2_) & (!i_6_) & (g14)) + ((!i_4_) & (i_5_) & (i_1_) & (i_2_) & (i_6_) & (g14)) + ((i_4_) & (i_5_) & (!i_1_) & (i_2_) & (i_6_) & (g14)));
	assign g461 = (((!i_3_) & (!i_6_) & (!i_8_) & (!g13)));
	assign g462 = (((!g27) & (!g28) & (!g36) & (!g461)) + ((!g27) & (!g28) & (g36) & (!g461)) + ((!g27) & (g28) & (g36) & (!g461)) + ((g27) & (!g28) & (!g36) & (!g461)) + ((g27) & (!g28) & (g36) & (!g461)) + ((g27) & (g28) & (!g36) & (!g461)) + ((g27) & (g28) & (g36) & (!g461)));
	assign g463 = (((!i_6_) & (!i_7_) & (!i_8_) & (!g71) & (g26)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g71) & (g26)) + ((!i_6_) & (!i_7_) & (i_8_) & (g71) & (!g26)) + ((!i_6_) & (!i_7_) & (i_8_) & (g71) & (g26)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g71) & (g26)) + ((!i_6_) & (i_7_) & (!i_8_) & (g71) & (g26)) + ((i_6_) & (i_7_) & (!i_8_) & (!g71) & (g26)) + ((i_6_) & (i_7_) & (!i_8_) & (g71) & (g26)));
	assign g464 = (((!g50) & (g47) & (!g94) & (g401)) + ((!g50) & (g47) & (g94) & (g401)) + ((g50) & (g47) & (!g94) & (g401)) + ((g50) & (g47) & (g94) & (!g401)) + ((g50) & (g47) & (g94) & (g401)));
	assign g465 = (((!g292) & (g327) & (!g363) & (!g463) & (!g464)));
	assign g466 = (((!g34) & (g323) & (!g460) & (g462) & (g465)));
	assign g467 = (((g154) & (g216) & (g445) & (g456) & (g459) & (g466)));
	assign g468 = (((!g8) & (!g45) & (!g13) & (!g165)) + ((!g8) & (!g45) & (g13) & (!g165)) + ((!g8) & (g45) & (!g13) & (!g165)) + ((!g8) & (g45) & (g13) & (!g165)) + ((g8) & (!g45) & (g13) & (!g165)) + ((g8) & (g45) & (!g13) & (!g165)) + ((g8) & (g45) & (g13) & (!g165)));
	assign g469 = (((!g21) & (!g6) & (!g23) & (!g24) & (!g3)) + ((!g21) & (!g6) & (!g23) & (!g24) & (g3)) + ((!g21) & (g6) & (!g23) & (!g24) & (!g3)) + ((!g21) & (g6) & (!g23) & (!g24) & (g3)) + ((!g21) & (g6) & (g23) & (!g24) & (g3)) + ((g21) & (g6) & (!g23) & (!g24) & (g3)) + ((g21) & (g6) & (g23) & (!g24) & (g3)));
	assign g470 = (((!g8) & (!g2) & (!g26) & (!g239) & (!g469)) + ((!g8) & (!g2) & (g26) & (!g239) & (!g469)) + ((!g8) & (g2) & (!g26) & (!g239) & (!g469)) + ((g8) & (!g2) & (!g26) & (!g239) & (!g469)) + ((g8) & (g2) & (!g26) & (!g239) & (!g469)));
	assign g471 = (((!g102) & (!g208) & (!g278) & (g40) & (g470)));
	assign g474 = (((!g42) & (!g38) & (g29) & (!g159)) + ((!g42) & (!g38) & (g29) & (g159)) + ((g42) & (!g38) & (!g29) & (g159)) + ((g42) & (!g38) & (g29) & (!g159)) + ((g42) & (!g38) & (g29) & (g159)) + ((g42) & (g38) & (!g29) & (g159)) + ((g42) & (g38) & (g29) & (g159)));
	assign g475 = (((g694) & (!g473) & (g400) & (!g409) & (!g474)));
	assign g477 = (((g50) & (i_6_) & (g63) & (g440)));
	assign g478 = (((!i_6_) & (i_7_) & (i_8_) & (g181) & (!g105) & (!g359)) + ((!i_6_) & (i_7_) & (i_8_) & (g181) & (!g105) & (g359)) + ((!i_6_) & (i_7_) & (i_8_) & (g181) & (g105) & (!g359)) + ((!i_6_) & (i_7_) & (i_8_) & (g181) & (g105) & (g359)) + ((i_6_) & (!i_7_) & (!i_8_) & (g181) & (!g105) & (!g359)) + ((i_6_) & (!i_7_) & (!i_8_) & (g181) & (!g105) & (g359)) + ((i_6_) & (!i_7_) & (!i_8_) & (g181) & (g105) & (!g359)) + ((i_6_) & (!i_7_) & (!i_8_) & (g181) & (g105) & (g359)) + ((i_6_) & (!i_7_) & (i_8_) & (!g181) & (!g105) & (!g359)) + ((i_6_) & (!i_7_) & (i_8_) & (!g181) & (!g105) & (g359)) + ((i_6_) & (!i_7_) & (i_8_) & (g181) & (!g105) & (!g359)) + ((i_6_) & (!i_7_) & (i_8_) & (g181) & (!g105) & (g359)) + ((i_6_) & (i_7_) & (!i_8_) & (!g181) & (!g105) & (g359)) + ((i_6_) & (i_7_) & (!i_8_) & (!g181) & (g105) & (g359)) + ((i_6_) & (i_7_) & (!i_8_) & (g181) & (!g105) & (g359)) + ((i_6_) & (i_7_) & (!i_8_) & (g181) & (g105) & (g359)));
	assign g479 = (((!g41) & (!g32) & (g343) & (g549) & (!g478)) + ((!g41) & (g32) & (g343) & (g549) & (!g478)) + ((g41) & (!g32) & (g343) & (g549) & (!g478)));
	assign g480 = (((!g43) & (!g92) & (g257) & (!g477) & (g479)));
	assign g481 = (((!g46) & (!g60) & (!g226) & (!g396) & (g456)) + ((!g46) & (g60) & (!g226) & (!g396) & (g456)) + ((g46) & (!g60) & (!g226) & (!g396) & (g456)));
	assign g483 = (((!g21) & (!g12) & (g6) & (!g13) & (g110)) + ((!g21) & (!g12) & (g6) & (g13) & (g110)) + ((!g21) & (g12) & (!g6) & (!g13) & (!g110)) + ((!g21) & (g12) & (!g6) & (!g13) & (g110)) + ((!g21) & (g12) & (g6) & (!g13) & (!g110)) + ((!g21) & (g12) & (g6) & (!g13) & (g110)) + ((!g21) & (g12) & (g6) & (g13) & (g110)));
	assign g484 = (((!g28) & (!g25) & (g12) & (g32) & (!g36)) + ((!g28) & (!g25) & (g12) & (g32) & (g36)) + ((g28) & (!g25) & (!g12) & (!g32) & (!g36)) + ((g28) & (!g25) & (!g12) & (g32) & (!g36)) + ((g28) & (!g25) & (g12) & (!g32) & (!g36)) + ((g28) & (!g25) & (g12) & (g32) & (!g36)) + ((g28) & (!g25) & (g12) & (g32) & (g36)));
	assign g485 = (((!g11) & (!g27) & (!g45) & (!g48) & (g2) & (!g24)) + ((!g11) & (!g27) & (!g45) & (!g48) & (g2) & (g24)) + ((!g11) & (!g27) & (!g45) & (g48) & (!g2) & (!g24)) + ((!g11) & (!g27) & (!g45) & (g48) & (g2) & (!g24)) + ((!g11) & (!g27) & (!g45) & (g48) & (g2) & (g24)) + ((!g11) & (!g27) & (g45) & (!g48) & (g2) & (!g24)) + ((!g11) & (!g27) & (g45) & (g48) & (g2) & (!g24)) + ((!g11) & (g27) & (!g45) & (!g48) & (g2) & (!g24)) + ((!g11) & (g27) & (!g45) & (g48) & (!g2) & (!g24)) + ((!g11) & (g27) & (!g45) & (g48) & (g2) & (!g24)) + ((!g11) & (g27) & (g45) & (!g48) & (g2) & (!g24)) + ((!g11) & (g27) & (g45) & (g48) & (g2) & (!g24)) + ((g11) & (!g27) & (!g45) & (!g48) & (g2) & (!g24)) + ((g11) & (!g27) & (!g45) & (!g48) & (g2) & (g24)) + ((g11) & (!g27) & (!g45) & (g48) & (!g2) & (!g24)) + ((g11) & (!g27) & (!g45) & (g48) & (g2) & (!g24)) + ((g11) & (!g27) & (!g45) & (g48) & (g2) & (g24)) + ((g11) & (g27) & (!g45) & (g48) & (!g2) & (!g24)) + ((g11) & (g27) & (!g45) & (g48) & (g2) & (!g24)));
	assign g486 = (((!g1) & (!g6) & (!g23) & (g3) & (!g49) & (!g110)) + ((!g1) & (!g6) & (!g23) & (g3) & (!g49) & (g110)) + ((!g1) & (!g6) & (!g23) & (g3) & (g49) & (!g110)) + ((!g1) & (!g6) & (!g23) & (g3) & (g49) & (g110)) + ((!g1) & (g6) & (!g23) & (!g3) & (g49) & (!g110)) + ((!g1) & (g6) & (!g23) & (!g3) & (g49) & (g110)) + ((!g1) & (g6) & (!g23) & (g3) & (!g49) & (!g110)) + ((!g1) & (g6) & (!g23) & (g3) & (!g49) & (g110)) + ((!g1) & (g6) & (!g23) & (g3) & (g49) & (!g110)) + ((!g1) & (g6) & (!g23) & (g3) & (g49) & (g110)) + ((!g1) & (g6) & (g23) & (!g3) & (g49) & (!g110)) + ((!g1) & (g6) & (g23) & (!g3) & (g49) & (g110)) + ((!g1) & (g6) & (g23) & (g3) & (!g49) & (g110)) + ((!g1) & (g6) & (g23) & (g3) & (g49) & (!g110)) + ((!g1) & (g6) & (g23) & (g3) & (g49) & (g110)) + ((g1) & (g6) & (!g23) & (!g3) & (g49) & (!g110)) + ((g1) & (g6) & (!g23) & (!g3) & (g49) & (g110)) + ((g1) & (g6) & (!g23) & (g3) & (!g49) & (g110)) + ((g1) & (g6) & (!g23) & (g3) & (g49) & (!g110)) + ((g1) & (g6) & (!g23) & (g3) & (g49) & (g110)) + ((g1) & (g6) & (g23) & (!g3) & (g49) & (!g110)) + ((g1) & (g6) & (g23) & (!g3) & (g49) & (g110)) + ((g1) & (g6) & (g23) & (g3) & (!g49) & (g110)) + ((g1) & (g6) & (g23) & (g3) & (g49) & (!g110)) + ((g1) & (g6) & (g23) & (g3) & (g49) & (g110)));
	assign g488 = (((!i_6_) & (!i_7_) & (!g188) & (!g129)) + ((!i_6_) & (!i_7_) & (!g188) & (g129)) + ((!i_6_) & (i_7_) & (!g188) & (!g129)) + ((!i_6_) & (i_7_) & (!g188) & (g129)) + ((i_6_) & (!i_7_) & (!g188) & (!g129)) + ((i_6_) & (i_7_) & (!g188) & (!g129)) + ((i_6_) & (i_7_) & (!g188) & (g129)));
	assign g489 = (((!i_6_) & (!g32) & (!g18) & (!g110) & (g488)) + ((!i_6_) & (!g32) & (!g18) & (g110) & (g488)) + ((!i_6_) & (g32) & (!g18) & (!g110) & (g488)) + ((!i_6_) & (g32) & (!g18) & (g110) & (g488)) + ((i_6_) & (!g32) & (!g18) & (!g110) & (g488)) + ((i_6_) & (!g32) & (!g18) & (g110) & (g488)) + ((i_6_) & (g32) & (!g18) & (!g110) & (g488)));
	assign g490 = (((g476) & (g482) & (g487) & (g489)));
	assign g492 = (((!g1) & (!g12) & (!g3) & (!g290)) + ((!g1) & (!g12) & (g3) & (!g290)) + ((!g1) & (g12) & (!g3) & (!g290)) + ((g1) & (!g12) & (!g3) & (!g290)) + ((g1) & (!g12) & (g3) & (!g290)) + ((g1) & (g12) & (!g3) & (!g290)) + ((g1) & (g12) & (g3) & (!g290)));
	assign g493 = (((!g11) & (!g41) & (!g45) & (!g29) & (!g141)) + ((!g11) & (!g41) & (g45) & (!g29) & (!g141)) + ((!g11) & (!g41) & (g45) & (g29) & (!g141)) + ((!g11) & (g41) & (g45) & (!g29) & (!g141)) + ((!g11) & (g41) & (g45) & (g29) & (!g141)) + ((g11) & (!g41) & (!g45) & (!g29) & (!g141)) + ((g11) & (!g41) & (!g45) & (!g29) & (g141)) + ((g11) & (!g41) & (g45) & (!g29) & (!g141)) + ((g11) & (!g41) & (g45) & (!g29) & (g141)) + ((g11) & (!g41) & (g45) & (g29) & (!g141)) + ((g11) & (!g41) & (g45) & (g29) & (g141)) + ((g11) & (g41) & (g45) & (!g29) & (!g141)) + ((g11) & (g41) & (g45) & (!g29) & (g141)) + ((g11) & (g41) & (g45) & (g29) & (!g141)) + ((g11) & (g41) & (g45) & (g29) & (g141)));
	assign g494 = (((!g21) & (!g48) & (!g49) & (!g110) & (!g364)) + ((!g21) & (!g48) & (!g49) & (g110) & (!g364)) + ((!g21) & (!g48) & (g49) & (!g110) & (!g364)) + ((!g21) & (!g48) & (g49) & (g110) & (!g364)) + ((!g21) & (g48) & (!g49) & (!g110) & (!g364)) + ((g21) & (!g48) & (!g49) & (!g110) & (!g364)) + ((g21) & (!g48) & (!g49) & (g110) & (!g364)) + ((g21) & (!g48) & (g49) & (!g110) & (!g364)) + ((g21) & (!g48) & (g49) & (g110) & (!g364)) + ((g21) & (g48) & (!g49) & (!g110) & (!g364)) + ((g21) & (g48) & (!g49) & (g110) & (!g364)));
	assign g495 = (((!g23) & (!g184) & (g492) & (g493) & (g494)) + ((g23) & (!g184) & (g492) & (g493) & (g494)) + ((g23) & (g184) & (g492) & (g493) & (g494)));
	assign g499 = (((!i_0_) & (!i_1_) & (!i_2_) & (!g194)) + ((!i_0_) & (!i_1_) & (!i_2_) & (g194)) + ((!i_0_) & (i_1_) & (!i_2_) & (g194)));
	assign g501 = (((!g23) & (!g71) & (!g294) & (!g88) & (!g212)) + ((g23) & (!g71) & (!g294) & (!g88) & (!g212)) + ((g23) & (!g71) & (!g294) & (g88) & (!g212)) + ((g23) & (g71) & (!g294) & (!g88) & (!g212)) + ((g23) & (g71) & (!g294) & (g88) & (!g212)));
	assign g502 = (((!g27) & (!g12) & (!g33) & (!g4) & (!g194)) + ((!g27) & (!g12) & (g33) & (!g4) & (!g194)) + ((!g27) & (g12) & (!g33) & (!g4) & (!g194)) + ((g27) & (!g12) & (!g33) & (!g4) & (!g194)) + ((g27) & (!g12) & (!g33) & (!g4) & (g194)) + ((g27) & (!g12) & (!g33) & (g4) & (!g194)) + ((g27) & (!g12) & (!g33) & (g4) & (g194)) + ((g27) & (!g12) & (g33) & (!g4) & (!g194)) + ((g27) & (!g12) & (g33) & (!g4) & (g194)) + ((g27) & (!g12) & (g33) & (g4) & (!g194)) + ((g27) & (!g12) & (g33) & (g4) & (g194)) + ((g27) & (g12) & (!g33) & (!g4) & (!g194)) + ((g27) & (g12) & (!g33) & (!g4) & (g194)) + ((g27) & (g12) & (!g33) & (g4) & (!g194)) + ((g27) & (g12) & (!g33) & (g4) & (g194)));
	assign g503 = (((!g174) & (!g277) & (g500) & (g501) & (g502)));
	assign g504 = (((!g6) & (!g59) & (!g88) & (g265)) + ((!g6) & (!g59) & (g88) & (g265)) + ((g6) & (!g59) & (!g88) & (g265)) + ((g6) & (!g59) & (g88) & (!g265)) + ((g6) & (!g59) & (g88) & (g265)) + ((g6) & (g59) & (g88) & (!g265)) + ((g6) & (g59) & (g88) & (g265)));
	assign g505 = (((!g37) & (!g129) & (g386) & (!g504)) + ((!g37) & (g129) & (g386) & (!g504)) + ((g37) & (!g129) & (g386) & (!g504)));
	assign g507 = (((g35) & (!g45) & (!g13)));
	assign g508 = (((!i_3_) & (!g50) & (!g127) & (g8) & (g84)) + ((!i_3_) & (!g50) & (g127) & (g8) & (g84)) + ((!i_3_) & (g50) & (!g127) & (g8) & (g84)) + ((!i_3_) & (g50) & (g127) & (g8) & (!g84)) + ((!i_3_) & (g50) & (g127) & (g8) & (g84)) + ((i_3_) & (!g50) & (!g127) & (g8) & (g84)) + ((i_3_) & (!g50) & (g127) & (g8) & (g84)) + ((i_3_) & (g50) & (!g127) & (g8) & (g84)) + ((i_3_) & (g50) & (g127) & (g8) & (g84)));
	assign g509 = (((!g63) & (!g6) & (!g129) & (!g507) & (!g508)) + ((!g63) & (!g6) & (g129) & (!g507) & (!g508)) + ((!g63) & (g6) & (!g129) & (!g507) & (!g508)) + ((g63) & (!g6) & (!g129) & (!g507) & (!g508)) + ((g63) & (g6) & (!g129) & (!g507) & (!g508)));
	assign g510 = (((g476) & (g496) & (g506) & (g509)));
	assign g511 = (((!g21) & (!g25) & (!g48) & (g2) & (!g13) & (!g38)) + ((!g21) & (!g25) & (!g48) & (g2) & (!g13) & (g38)) + ((!g21) & (!g25) & (!g48) & (g2) & (g13) & (!g38)) + ((!g21) & (!g25) & (g48) & (!g2) & (!g13) & (!g38)) + ((!g21) & (!g25) & (g48) & (!g2) & (!g13) & (g38)) + ((!g21) & (!g25) & (g48) & (!g2) & (g13) & (!g38)) + ((!g21) & (!g25) & (g48) & (!g2) & (g13) & (g38)) + ((!g21) & (!g25) & (g48) & (g2) & (!g13) & (!g38)) + ((!g21) & (!g25) & (g48) & (g2) & (!g13) & (g38)) + ((!g21) & (!g25) & (g48) & (g2) & (g13) & (!g38)) + ((!g21) & (!g25) & (g48) & (g2) & (g13) & (g38)) + ((!g21) & (g25) & (!g48) & (g2) & (!g13) & (!g38)) + ((!g21) & (g25) & (!g48) & (g2) & (!g13) & (g38)) + ((!g21) & (g25) & (g48) & (g2) & (!g13) & (!g38)) + ((!g21) & (g25) & (g48) & (g2) & (!g13) & (g38)) + ((g21) & (!g25) & (!g48) & (g2) & (!g13) & (!g38)) + ((g21) & (!g25) & (!g48) & (g2) & (g13) & (!g38)) + ((g21) & (!g25) & (g48) & (g2) & (!g13) & (!g38)) + ((g21) & (!g25) & (g48) & (g2) & (g13) & (!g38)));
	assign g512 = (((!g42) & (!g12) & (!g59) & (g7)) + ((!g42) & (g12) & (!g59) & (g7)) + ((g42) & (!g12) & (!g59) & (g7)) + ((g42) & (g12) & (!g59) & (!g7)) + ((g42) & (g12) & (!g59) & (g7)));
	assign g513 = (((!g27) & (!g45) & (g23) & (!g512)) + ((!g27) & (g45) & (!g23) & (!g512)) + ((!g27) & (g45) & (g23) & (!g512)) + ((g27) & (!g45) & (!g23) & (!g512)) + ((g27) & (!g45) & (g23) & (!g512)) + ((g27) & (g45) & (!g23) & (!g512)) + ((g27) & (g45) & (g23) & (!g512)));
	assign g514 = (((!g41) & (!g21) & (!g3) & (!g29) & (!g265)) + ((!g41) & (!g21) & (!g3) & (g29) & (!g265)) + ((!g41) & (!g21) & (g3) & (!g29) & (!g265)) + ((!g41) & (g21) & (!g3) & (!g29) & (!g265)) + ((!g41) & (g21) & (!g3) & (!g29) & (g265)) + ((!g41) & (g21) & (!g3) & (g29) & (!g265)) + ((!g41) & (g21) & (!g3) & (g29) & (g265)) + ((!g41) & (g21) & (g3) & (!g29) & (!g265)) + ((g41) & (!g21) & (!g3) & (!g29) & (!g265)) + ((g41) & (!g21) & (!g3) & (g29) & (!g265)) + ((g41) & (g21) & (!g3) & (!g29) & (!g265)) + ((g41) & (g21) & (!g3) & (!g29) & (g265)) + ((g41) & (g21) & (!g3) & (g29) & (!g265)) + ((g41) & (g21) & (!g3) & (g29) & (g265)));
	assign g515 = (((!g134) & (!g413) & (!g457) & (!g472) & (g514)) + ((!g134) & (!g413) & (!g457) & (g472) & (g514)) + ((g134) & (!g413) & (!g457) & (!g472) & (g514)));
	assign g516 = (((!g28) & (g32) & (g67) & (!g181)) + ((!g28) & (g32) & (g67) & (g181)) + ((g28) & (!g32) & (!g67) & (g181)) + ((g28) & (!g32) & (g67) & (g181)) + ((g28) & (g32) & (!g67) & (g181)) + ((g28) & (g32) & (g67) & (!g181)) + ((g28) & (g32) & (g67) & (g181)));
	assign g517 = (((!g314) & (!g293) & (g236) & (!g516)));
	assign g519 = (((!g13) & (!g123) & (!g387) & (!g458)) + ((g13) & (!g123) & (!g387) & (!g458)) + ((g13) & (g123) & (!g387) & (!g458)));
	assign g520 = (((!g431) & (g487) & (g506) & (g518) & (g519)));
	assign g521 = (((!g8) & (!g117) & (!g428)) + ((!g8) & (g117) & (!g428)) + ((g8) & (!g117) & (!g428)));
	assign g522 = (((!i_4_) & (!i_5_) & (!g63) & (!g65) & (!g472) & (g521)) + ((!i_4_) & (!i_5_) & (!g63) & (!g65) & (g472) & (g521)) + ((!i_4_) & (!i_5_) & (!g63) & (g65) & (!g472) & (g521)) + ((!i_4_) & (!i_5_) & (!g63) & (g65) & (g472) & (g521)) + ((!i_4_) & (!i_5_) & (g63) & (!g65) & (!g472) & (g521)) + ((!i_4_) & (i_5_) & (!g63) & (!g65) & (!g472) & (g521)) + ((!i_4_) & (i_5_) & (!g63) & (!g65) & (g472) & (g521)) + ((!i_4_) & (i_5_) & (!g63) & (g65) & (!g472) & (g521)) + ((!i_4_) & (i_5_) & (!g63) & (g65) & (g472) & (g521)) + ((!i_4_) & (i_5_) & (g63) & (!g65) & (!g472) & (g521)) + ((!i_4_) & (i_5_) & (g63) & (!g65) & (g472) & (g521)) + ((i_4_) & (!i_5_) & (!g63) & (!g65) & (!g472) & (g521)) + ((i_4_) & (!i_5_) & (!g63) & (!g65) & (g472) & (g521)) + ((i_4_) & (!i_5_) & (!g63) & (g65) & (!g472) & (g521)) + ((i_4_) & (!i_5_) & (!g63) & (g65) & (g472) & (g521)) + ((i_4_) & (!i_5_) & (g63) & (!g65) & (!g472) & (g521)) + ((i_4_) & (!i_5_) & (g63) & (!g65) & (g472) & (g521)) + ((i_4_) & (i_5_) & (!g63) & (!g65) & (!g472) & (g521)) + ((i_4_) & (i_5_) & (!g63) & (!g65) & (g472) & (g521)) + ((i_4_) & (i_5_) & (!g63) & (g65) & (!g472) & (g521)) + ((i_4_) & (i_5_) & (!g63) & (g65) & (g472) & (g521)) + ((i_4_) & (i_5_) & (g63) & (!g65) & (!g472) & (g521)) + ((i_4_) & (i_5_) & (g63) & (!g65) & (g472) & (g521)));
	assign g523 = (((g482) & (g496) & (g518) & (g522)));
	assign g525 = (((i_6_) & (!i_7_) & (!i_8_) & (!g45) & (!g3) & (g110)) + ((i_6_) & (!i_7_) & (!i_8_) & (!g45) & (g3) & (g110)) + ((i_6_) & (!i_7_) & (i_8_) & (!g45) & (!g3) & (g110)) + ((i_6_) & (!i_7_) & (i_8_) & (!g45) & (g3) & (g110)) + ((i_6_) & (i_7_) & (!i_8_) & (!g45) & (!g3) & (g110)) + ((i_6_) & (i_7_) & (!i_8_) & (!g45) & (g3) & (g110)) + ((i_6_) & (i_7_) & (!i_8_) & (g45) & (g3) & (g110)) + ((i_6_) & (i_7_) & (i_8_) & (!g45) & (!g3) & (g110)) + ((i_6_) & (i_7_) & (i_8_) & (!g45) & (g3) & (g110)));
	assign g526 = (((!i_6_) & (i_7_) & (!i_8_) & (!g21) & (!g25) & (!g110)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g21) & (!g25) & (g110)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g21) & (g25) & (g110)) + ((!i_6_) & (i_7_) & (i_8_) & (!g21) & (!g25) & (!g110)) + ((!i_6_) & (i_7_) & (i_8_) & (!g21) & (!g25) & (g110)) + ((i_6_) & (i_7_) & (!i_8_) & (!g21) & (!g25) & (!g110)) + ((i_6_) & (i_7_) & (!i_8_) & (!g21) & (!g25) & (g110)) + ((i_6_) & (i_7_) & (i_8_) & (!g21) & (!g25) & (!g110)) + ((i_6_) & (i_7_) & (i_8_) & (!g21) & (!g25) & (g110)));
	assign g527 = (((!i_6_) & (!i_7_) & (!i_8_) & (!g46) & (g184)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g46) & (!g184)) + ((!i_6_) & (!i_7_) & (!i_8_) & (g46) & (g184)) + ((!i_6_) & (!i_7_) & (i_8_) & (!g46) & (g184)) + ((!i_6_) & (!i_7_) & (i_8_) & (g46) & (g184)) + ((!i_6_) & (i_7_) & (!i_8_) & (!g46) & (g184)) + ((!i_6_) & (i_7_) & (!i_8_) & (g46) & (g184)));
	assign g529 = (((!i_6_) & (i_7_) & (!i_8_) & (g189) & (!g161)) + ((!i_6_) & (i_7_) & (!i_8_) & (g189) & (g161)) + ((!i_6_) & (i_7_) & (i_8_) & (g189) & (!g161)) + ((!i_6_) & (i_7_) & (i_8_) & (g189) & (g161)) + ((i_6_) & (!i_7_) & (i_8_) & (!g189) & (g161)) + ((i_6_) & (!i_7_) & (i_8_) & (g189) & (!g161)) + ((i_6_) & (!i_7_) & (i_8_) & (g189) & (g161)) + ((i_6_) & (i_7_) & (!i_8_) & (!g189) & (g161)) + ((i_6_) & (i_7_) & (!i_8_) & (g189) & (g161)) + ((i_6_) & (i_7_) & (i_8_) & (!g189) & (g161)) + ((i_6_) & (i_7_) & (i_8_) & (g189) & (g161)));
	assign g530 = (((!g25) & (!g23) & (g38) & (!g491)) + ((!g25) & (g23) & (!g38) & (!g491)) + ((!g25) & (g23) & (g38) & (!g491)) + ((g25) & (!g23) & (!g38) & (!g491)) + ((g25) & (!g23) & (g38) & (!g491)) + ((g25) & (g23) & (!g38) & (!g491)) + ((g25) & (g23) & (g38) & (!g491)));
	assign g532 = (((!g524) & (g528) & (g531)));
	assign g534 = (((!i_0_) & (!i_1_) & (!i_2_) & (!g2) & (!g59)) + ((!i_0_) & (!i_1_) & (!i_2_) & (!g2) & (g59)) + ((!i_0_) & (!i_1_) & (!i_2_) & (g2) & (!g59)) + ((!i_0_) & (!i_1_) & (!i_2_) & (g2) & (g59)) + ((!i_0_) & (i_1_) & (!i_2_) & (g2) & (!g59)));
	assign g535 = (((!g6) & (!g23) & (g189) & (!g99)) + ((!g6) & (!g23) & (g189) & (g99)) + ((g6) & (!g23) & (!g189) & (g99)) + ((g6) & (!g23) & (g189) & (!g99)) + ((g6) & (!g23) & (g189) & (g99)) + ((g6) & (g23) & (!g189) & (g99)) + ((g6) & (g23) & (g189) & (g99)));
	assign g537 = (((!g533) & (g531) & (g536)));
	assign g539 = (((!i_4_) & (!i_6_) & (!g6) & (!g161) & (g472)) + ((!i_4_) & (!i_6_) & (!g6) & (g161) & (g472)) + ((!i_4_) & (!i_6_) & (g6) & (!g161) & (g472)) + ((!i_4_) & (!i_6_) & (g6) & (g161) & (!g472)) + ((!i_4_) & (!i_6_) & (g6) & (g161) & (g472)) + ((!i_4_) & (i_6_) & (g6) & (g161) & (!g472)) + ((!i_4_) & (i_6_) & (g6) & (g161) & (g472)) + ((i_4_) & (!i_6_) & (g6) & (g161) & (!g472)) + ((i_4_) & (!i_6_) & (g6) & (g161) & (g472)) + ((i_4_) & (i_6_) & (g6) & (g161) & (!g472)) + ((i_4_) & (i_6_) & (g6) & (g161) & (g472)));
	assign g540 = (((!g497) & (!g524) & (!g538) & (g536) & (!g539)));
	assign g541 = (((!i_4_) & (!i_5_) & (!i_6_) & (!g63) & (g472)) + ((!i_4_) & (!i_5_) & (!i_6_) & (g63) & (g472)) + ((!i_4_) & (!i_5_) & (i_6_) & (g63) & (g472)));
	assign g542 = (((!g533) & (!g538) & (!g541) & (g528)));
	assign g543 = (((g515) & (g544)));
	assign g544 = (((!g545) & (g546)) + ((g545) & (!g546)) + ((g545) & (g546)));
	assign g545 = (((!i_6_) & (g547)));
	assign g546 = (((i_6_) & (g548)));
	assign g547 = (((!i_8_) & (!g88) & (!i_7_)) + ((!i_8_) & (!g88) & (i_7_)) + ((!i_8_) & (g88) & (!i_7_)) + ((i_8_) & (!g88) & (!i_7_)) + ((i_8_) & (!g88) & (i_7_)) + ((i_8_) & (g88) & (i_7_)));
	assign g548 = (((!g98) & (!i_8_) & (!g73) & (!i_7_)) + ((!g98) & (!i_8_) & (!g73) & (i_7_)) + ((!g98) & (!i_8_) & (g73) & (!i_7_)) + ((!g98) & (i_8_) & (!g73) & (!i_7_)) + ((!g98) & (i_8_) & (!g73) & (i_7_)) + ((!g98) & (i_8_) & (g73) & (!i_7_)) + ((!g98) & (i_8_) & (g73) & (i_7_)) + ((g98) & (!i_8_) & (!g73) & (!i_7_)) + ((g98) & (!i_8_) & (g73) & (!i_7_)) + ((g98) & (i_8_) & (!g73) & (!i_7_)) + ((g98) & (i_8_) & (!g73) & (i_7_)) + ((g98) & (i_8_) & (g73) & (!i_7_)) + ((g98) & (i_8_) & (g73) & (i_7_)));
	assign g549 = (((!g550) & (g551)) + ((g550) & (!g551)) + ((g550) & (g551)));
	assign g550 = (((!i_0_) & (g552)));
	assign g551 = (((i_0_) & (g554)));
	assign g552 = (((!i_1_) & (g553)) + ((i_1_) & (!g553)) + ((i_1_) & (g553)));
	assign g553 = (((!i_1_) & (i_2_)));
	assign g554 = (((!g555) & (g556)) + ((g555) & (!g556)) + ((g555) & (g556)));
	assign g555 = (((!i_1_) & (g557)));
	assign g556 = (((i_1_) & (g558)));
	assign g557 = (((!g36) & (!g23) & (!g6) & (i_2_)) + ((!g36) & (!g23) & (g6) & (i_2_)) + ((!g36) & (g23) & (!g6) & (!i_2_)) + ((!g36) & (g23) & (!g6) & (i_2_)) + ((!g36) & (g23) & (g6) & (i_2_)) + ((g36) & (!g23) & (!g6) & (!i_2_)) + ((g36) & (!g23) & (!g6) & (i_2_)) + ((g36) & (!g23) & (g6) & (!i_2_)) + ((g36) & (!g23) & (g6) & (i_2_)) + ((g36) & (g23) & (!g6) & (!i_2_)) + ((g36) & (g23) & (!g6) & (i_2_)) + ((g36) & (g23) & (g6) & (!i_2_)) + ((g36) & (g23) & (g6) & (i_2_)));
	assign g558 = (((!g16) & (!i_2_)) + ((!g16) & (i_2_)) + ((g16) & (i_2_)));
	assign g559 = (((!g560) & (g561)) + ((g560) & (!g561)) + ((g560) & (g561)));
	assign g560 = (((!g243) & (g562)));
	assign g561 = (((g243) & (g565)));
	assign g562 = (((!g563) & (g564)) + ((g563) & (!g564)) + ((g563) & (g564)));
	assign g563 = (((!i_8_) & (g568)));
	assign g564 = (((i_8_) & (g569)));
	assign g565 = (((!g566) & (g567)) + ((g566) & (!g567)) + ((g566) & (g567)));
	assign g566 = (((!i_8_) & (g570)));
	assign g567 = (((i_8_) & (g571)));
	assign g568 = (((g448) & (g449) & (g447)));
	assign g569 = (((g448) & (g449) & (g447)));
	assign g570 = (((g448) & (g449) & (i_7_) & (g447)));
	assign g571 = (((g448) & (g449) & (i_6_) & (g447)));
	assign g572 = (((!g573) & (g574)) + ((g573) & (!g574)) + ((g573) & (g574)));
	assign g573 = (((!i_6_) & (g575)));
	assign g574 = (((i_6_) & (g578)));
	assign g575 = (((!g576) & (g577)) + ((g576) & (!g577)) + ((g576) & (g577)));
	assign g576 = (((!i_8_) & (g580)));
	assign g577 = (((i_8_) & (g581)));
	assign g578 = (((!i_8_) & (g579)) + ((i_8_) & (!g579)) + ((i_8_) & (g579)));
	assign g579 = (((!i_8_) & (g582)));
	assign g580 = (((!g59) & (!g25) & (i_7_)) + ((!g59) & (g25) & (!i_7_)) + ((!g59) & (g25) & (i_7_)) + ((g59) & (!g25) & (!i_7_)) + ((g59) & (!g25) & (i_7_)) + ((g59) & (g25) & (!i_7_)) + ((g59) & (g25) & (i_7_)));
	assign g581 = (((!g59) & (g13)) + ((g59) & (!g13)) + ((g59) & (g13)));
	assign g582 = (((!i_7_) & (g105)) + ((i_7_) & (!g105)) + ((i_7_) & (g105)));
	assign g583 = (((!g584) & (g585)) + ((g584) & (!g585)) + ((g584) & (g585)));
	assign g584 = (((!g359) & (g586)));
	assign g585 = (((g359) & (g589)));
	assign g586 = (((!g587) & (g588)) + ((g587) & (!g588)) + ((g587) & (g588)));
	assign g587 = (((!i_6_) & (g592)));
	assign g588 = (((i_6_) & (g593)));
	assign g589 = (((!g590) & (g591)) + ((g590) & (!g591)) + ((g590) & (g591)));
	assign g590 = (((!i_6_) & (g594)));
	assign g591 = (((i_6_) & (g595)));
	assign g592 = (((!i_8_) & (!i_7_) & (!g105) & (g392)) + ((!i_8_) & (!i_7_) & (g105) & (g392)) + ((!i_8_) & (i_7_) & (g105) & (g392)) + ((i_8_) & (!i_7_) & (!g105) & (g392)) + ((i_8_) & (!i_7_) & (g105) & (g392)) + ((i_8_) & (i_7_) & (!g105) & (g392)) + ((i_8_) & (i_7_) & (g105) & (g392)));
	assign g593 = (((!i_8_) & (!i_7_) & (!g98) & (g392)) + ((!i_8_) & (i_7_) & (!g98) & (g392)) + ((i_8_) & (!i_7_) & (!g98) & (g392)) + ((i_8_) & (!i_7_) & (g98) & (g392)) + ((i_8_) & (i_7_) & (!g98) & (g392)));
	assign g594 = (((!i_8_) & (!i_7_) & (g392)) + ((i_8_) & (!i_7_) & (g392)) + ((i_8_) & (i_7_) & (g392)));
	assign g595 = (((!i_8_) & (!i_7_) & (!g98) & (g392)) + ((!i_8_) & (i_7_) & (!g98) & (g392)) + ((i_8_) & (!i_7_) & (!g98) & (g392)) + ((i_8_) & (!i_7_) & (g98) & (g392)) + ((i_8_) & (i_7_) & (!g98) & (g392)));
	assign g596 = (((!g597) & (g598)) + ((g597) & (!g598)) + ((g597) & (g598)));
	assign g597 = (((!i_6_) & (g599)));
	assign g598 = (((i_6_) & (g601)));
	assign g599 = (((!i_7_) & (g600)) + ((i_7_) & (!g600)) + ((i_7_) & (g600)));
	assign g600 = (((!i_7_) & (g604)));
	assign g601 = (((!g602) & (g603)) + ((g602) & (!g603)) + ((g602) & (g603)));
	assign g602 = (((!i_7_) & (g605)));
	assign g603 = (((i_7_) & (g606)));
	assign g604 = (((!g59) & (!g25) & (!i_8_)) + ((!g59) & (g25) & (!i_8_)) + ((!g59) & (g25) & (i_8_)) + ((g59) & (!g25) & (!i_8_)) + ((g59) & (!g25) & (i_8_)) + ((g59) & (g25) & (!i_8_)) + ((g59) & (g25) & (i_8_)));
	assign g605 = (((!g98) & (!i_8_)) + ((!g98) & (i_8_)) + ((g98) & (!i_8_)));
	assign g606 = (((!g25) & (g21)) + ((g25) & (!g21)) + ((g25) & (g21)));
	assign g607 = (((!g608) & (g609)) + ((g608) & (!g609)) + ((g608) & (g609)));
	assign g608 = (((!g6) & (g610)));
	assign g609 = (((g6) & (g612)));
	assign g610 = (((!g11) & (g611)) + ((g11) & (!g611)) + ((g11) & (g611)));
	assign g611 = (((!g11) & (g615)));
	assign g612 = (((!g613) & (g614)) + ((g613) & (!g614)) + ((g613) & (g614)));
	assign g613 = (((!g11) & (g616)));
	assign g614 = (((g11) & (g617)));
	assign g615 = (((!g13) & (!g47)) + ((g13) & (!g47)) + ((g13) & (g47)));
	assign g616 = (((!g13) & (g24) & (!g47) & (!g99)) + ((g13) & (g24) & (!g47) & (!g99)) + ((g13) & (g24) & (g47) & (!g99)));
	assign g617 = (((!g24) & (g36) & (!g99)) + ((g24) & (!g36) & (!g99)) + ((g24) & (g36) & (!g99)));
	assign g619 = (((!g11) & (g621)));
	assign g620 = (((g11) & (g624)));
	assign g621 = (((!g622) & (g623)) + ((g622) & (!g623)) + ((g622) & (g623)));
	assign g622 = (((!i_8_) & (g627)));
	assign g623 = (((i_8_) & (g628)));
	assign g624 = (((!g625) & (g626)) + ((g625) & (!g626)) + ((g625) & (g626)));
	assign g625 = (((!i_8_) & (g629)));
	assign g626 = (((i_8_) & (g630)));
	assign g627 = (((!i_6_) & (!g46)) + ((!i_6_) & (g46)) + ((i_6_) & (!g46)));
	assign g628 = (((!g77) & (!i_6_) & (!i_7_) & (!g1)) + ((!g77) & (!i_6_) & (!i_7_) & (g1)) + ((!g77) & (!i_6_) & (i_7_) & (!g1)) + ((!g77) & (!i_6_) & (i_7_) & (g1)) + ((!g77) & (i_6_) & (!i_7_) & (g1)) + ((!g77) & (i_6_) & (i_7_) & (!g1)) + ((!g77) & (i_6_) & (i_7_) & (g1)) + ((g77) & (!i_6_) & (i_7_) & (!g1)) + ((g77) & (!i_6_) & (i_7_) & (g1)) + ((g77) & (i_6_) & (!i_7_) & (g1)) + ((g77) & (i_6_) & (i_7_) & (!g1)) + ((g77) & (i_6_) & (i_7_) & (g1)));
	assign g629 = (((!i_6_) & (!g46)) + ((!i_6_) & (g46)) + ((i_6_) & (!g46)));
	assign g630 = (((!g77) & (!i_6_) & (!i_7_)) + ((!g77) & (!i_6_) & (i_7_)) + ((!g77) & (i_6_) & (!i_7_)) + ((!g77) & (i_6_) & (i_7_)) + ((g77) & (!i_6_) & (i_7_)) + ((g77) & (i_6_) & (!i_7_)) + ((g77) & (i_6_) & (i_7_)));
	assign g632 = (((!g35) & (g634)));
	assign g633 = (((g35) & (g637)));
	assign g634 = (((!g635) & (g636)) + ((g635) & (!g636)) + ((g635) & (g636)));
	assign g635 = (((!i_5_) & (g640)));
	assign g636 = (((i_5_) & (g641)));
	assign g637 = (((!g638) & (g639)) + ((g638) & (!g639)) + ((g638) & (g639)));
	assign g638 = (((!i_5_) & (g642)));
	assign g639 = (((i_5_) & (g643)));
	assign g640 = (((!i_4_) & (!g121)) + ((!i_4_) & (g121)) + ((i_4_) & (!g121)));
	assign g641 = (((!g95) & (!i_4_) & (!i_6_)) + ((!g95) & (!i_4_) & (i_6_)) + ((!g95) & (i_4_) & (!i_6_)) + ((!g95) & (i_4_) & (i_6_)) + ((g95) & (!i_4_) & (!i_6_)) + ((g95) & (!i_4_) & (i_6_)) + ((g95) & (i_4_) & (i_6_)));
	assign g642 = (((!i_4_) & (!g121)) + ((!i_4_) & (g121)) + ((i_4_) & (!g121)));
	assign g643 = (((!g95) & (!i_4_) & (!i_6_) & (!g42)) + ((!g95) & (!i_4_) & (i_6_) & (!g42)) + ((!g95) & (i_4_) & (!i_6_) & (!g42)) + ((!g95) & (i_4_) & (!i_6_) & (g42)) + ((!g95) & (i_4_) & (i_6_) & (!g42)) + ((!g95) & (i_4_) & (i_6_) & (g42)) + ((g95) & (!i_4_) & (!i_6_) & (!g42)) + ((g95) & (!i_4_) & (i_6_) & (!g42)) + ((g95) & (i_4_) & (i_6_) & (!g42)) + ((g95) & (i_4_) & (i_6_) & (g42)));
	assign g644 = (((!g645) & (g646)) + ((g645) & (!g646)) + ((g645) & (g646)));
	assign g645 = (((!g42) & (g647)));
	assign g646 = (((g42) & (g650)));
	assign g647 = (((!g648) & (g649)) + ((g648) & (!g649)) + ((g648) & (g649)));
	assign g648 = (((!i_6_) & (g653)));
	assign g649 = (((i_6_) & (g654)));
	assign g650 = (((!g651) & (g652)) + ((g651) & (!g652)) + ((g651) & (g652)));
	assign g651 = (((!i_6_) & (g655)));
	assign g652 = (((i_6_) & (g656)));
	assign g653 = (((!g24) & (!i_8_) & (!g36) & (i_7_)) + ((!g24) & (!i_8_) & (g36) & (!i_7_)) + ((!g24) & (!i_8_) & (g36) & (i_7_)) + ((!g24) & (i_8_) & (!g36) & (!i_7_)) + ((!g24) & (i_8_) & (!g36) & (i_7_)) + ((!g24) & (i_8_) & (g36) & (!i_7_)) + ((!g24) & (i_8_) & (g36) & (i_7_)) + ((g24) & (!i_8_) & (!g36) & (!i_7_)) + ((g24) & (!i_8_) & (!g36) & (i_7_)) + ((g24) & (!i_8_) & (g36) & (!i_7_)) + ((g24) & (!i_8_) & (g36) & (i_7_)) + ((g24) & (i_8_) & (!g36) & (!i_7_)) + ((g24) & (i_8_) & (!g36) & (i_7_)) + ((g24) & (i_8_) & (g36) & (!i_7_)) + ((g24) & (i_8_) & (g36) & (i_7_)));
	assign g654 = (((!g24) & (!i_8_) & (!g45) & (!i_7_)) + ((!g24) & (!i_8_) & (!g45) & (i_7_)) + ((!g24) & (!i_8_) & (g45) & (!i_7_)) + ((!g24) & (!i_8_) & (g45) & (i_7_)) + ((!g24) & (i_8_) & (!g45) & (i_7_)) + ((!g24) & (i_8_) & (g45) & (!i_7_)) + ((!g24) & (i_8_) & (g45) & (i_7_)) + ((g24) & (!i_8_) & (!g45) & (!i_7_)) + ((g24) & (!i_8_) & (!g45) & (i_7_)) + ((g24) & (!i_8_) & (g45) & (!i_7_)) + ((g24) & (!i_8_) & (g45) & (i_7_)) + ((g24) & (i_8_) & (!g45) & (!i_7_)) + ((g24) & (i_8_) & (!g45) & (i_7_)) + ((g24) & (i_8_) & (g45) & (!i_7_)) + ((g24) & (i_8_) & (g45) & (i_7_)));
	assign g655 = (((!g24) & (!i_8_) & (!g36) & (i_7_)) + ((!g24) & (!i_8_) & (g36) & (!i_7_)) + ((!g24) & (!i_8_) & (g36) & (i_7_)) + ((!g24) & (i_8_) & (!g36) & (!i_7_)) + ((!g24) & (i_8_) & (!g36) & (i_7_)) + ((!g24) & (i_8_) & (g36) & (!i_7_)) + ((!g24) & (i_8_) & (g36) & (i_7_)) + ((g24) & (!i_8_) & (!g36) & (!i_7_)) + ((g24) & (!i_8_) & (!g36) & (i_7_)) + ((g24) & (!i_8_) & (g36) & (!i_7_)) + ((g24) & (!i_8_) & (g36) & (i_7_)) + ((g24) & (i_8_) & (!g36) & (!i_7_)) + ((g24) & (i_8_) & (!g36) & (i_7_)) + ((g24) & (i_8_) & (g36) & (!i_7_)) + ((g24) & (i_8_) & (g36) & (i_7_)));
	assign g656 = (((!g24) & (!i_8_) & (!g45) & (i_7_)) + ((!g24) & (!i_8_) & (g45) & (!i_7_)) + ((!g24) & (!i_8_) & (g45) & (i_7_)) + ((!g24) & (i_8_) & (!g45) & (i_7_)) + ((!g24) & (i_8_) & (g45) & (!i_7_)) + ((!g24) & (i_8_) & (g45) & (i_7_)) + ((g24) & (!i_8_) & (!g45) & (i_7_)) + ((g24) & (!i_8_) & (g45) & (!i_7_)) + ((g24) & (!i_8_) & (g45) & (i_7_)) + ((g24) & (i_8_) & (!g45) & (!i_7_)) + ((g24) & (i_8_) & (!g45) & (i_7_)) + ((g24) & (i_8_) & (g45) & (!i_7_)) + ((g24) & (i_8_) & (g45) & (i_7_)));
	assign g657 = (((!g658) & (g659)) + ((g658) & (!g659)) + ((g658) & (g659)));
	assign g658 = (((!g23) & (g660)));
	assign g659 = (((g23) & (g663)));
	assign g660 = (((!g661) & (g662)) + ((g661) & (!g662)) + ((g661) & (g662)));
	assign g661 = (((!i_2_) & (g666)));
	assign g662 = (((i_2_) & (g667)));
	assign g663 = (((!g664) & (g665)) + ((g664) & (!g665)) + ((g664) & (g665)));
	assign g664 = (((!i_2_) & (g668)));
	assign g665 = (((i_2_) & (g669)));
	assign g666 = (((!i_0_) & (!g187) & (!i_1_) & (!g38)) + ((!i_0_) & (!g187) & (!i_1_) & (g38)) + ((!i_0_) & (!g187) & (i_1_) & (!g38)) + ((!i_0_) & (!g187) & (i_1_) & (g38)) + ((!i_0_) & (g187) & (!i_1_) & (!g38)) + ((!i_0_) & (g187) & (!i_1_) & (g38)) + ((!i_0_) & (g187) & (i_1_) & (!g38)) + ((!i_0_) & (g187) & (i_1_) & (g38)) + ((i_0_) & (!g187) & (i_1_) & (!g38)) + ((i_0_) & (!g187) & (i_1_) & (g38)) + ((i_0_) & (g187) & (!i_1_) & (g38)) + ((i_0_) & (g187) & (i_1_) & (!g38)) + ((i_0_) & (g187) & (i_1_) & (g38)));
	assign g667 = (((!i_0_) & (!i_7_) & (!g38)) + ((!i_0_) & (!i_7_) & (g38)) + ((!i_0_) & (i_7_) & (!g38)) + ((!i_0_) & (i_7_) & (g38)) + ((i_0_) & (!i_7_) & (!g38)) + ((i_0_) & (!i_7_) & (g38)) + ((i_0_) & (i_7_) & (g38)));
	assign g668 = (((!i_0_) & (!g187) & (!i_1_)) + ((!i_0_) & (!g187) & (i_1_)) + ((!i_0_) & (g187) & (!i_1_)) + ((!i_0_) & (g187) & (i_1_)) + ((i_0_) & (!g187) & (i_1_)) + ((i_0_) & (g187) & (!i_1_)) + ((i_0_) & (g187) & (i_1_)));
	assign g669 = (((!i_0_) & (!i_7_) & (!g38)) + ((!i_0_) & (!i_7_) & (g38)) + ((!i_0_) & (i_7_) & (!g38)) + ((!i_0_) & (i_7_) & (g38)) + ((i_0_) & (!i_7_) & (!g38)) + ((i_0_) & (!i_7_) & (g38)) + ((i_0_) & (i_7_) & (g38)));
	assign g671 = (((!g41) & (g673)));
	assign g672 = (((g41) & (g676)));
	assign g673 = (((!g674) & (g675)) + ((g674) & (!g675)) + ((g674) & (g675)));
	assign g674 = (((!i_4_) & (g679)));
	assign g675 = (((i_4_) & (g680)));
	assign g676 = (((!g677) & (g678)) + ((g677) & (!g678)) + ((g677) & (g678)));
	assign g677 = (((!i_4_) & (g681)));
	assign g678 = (((i_4_) & (g682)));
	assign g679 = (((!g1) & (!i_5_) & (!g12) & (!i_3_)) + ((!g1) & (!i_5_) & (!g12) & (i_3_)) + ((!g1) & (!i_5_) & (g12) & (!i_3_)) + ((!g1) & (i_5_) & (!g12) & (!i_3_)) + ((!g1) & (i_5_) & (!g12) & (i_3_)) + ((!g1) & (i_5_) & (g12) & (!i_3_)) + ((!g1) & (i_5_) & (g12) & (i_3_)) + ((g1) & (!i_5_) & (!g12) & (!i_3_)) + ((g1) & (!i_5_) & (!g12) & (i_3_)) + ((g1) & (!i_5_) & (g12) & (!i_3_)) + ((g1) & (!i_5_) & (g12) & (i_3_)) + ((g1) & (i_5_) & (!g12) & (!i_3_)) + ((g1) & (i_5_) & (!g12) & (i_3_)) + ((g1) & (i_5_) & (g12) & (!i_3_)) + ((g1) & (i_5_) & (g12) & (i_3_)));
	assign g680 = (((!g1) & (!i_5_) & (!g28) & (!i_3_)) + ((!g1) & (!i_5_) & (!g28) & (i_3_)) + ((!g1) & (!i_5_) & (g28) & (!i_3_)) + ((!g1) & (i_5_) & (!g28) & (!i_3_)) + ((!g1) & (i_5_) & (!g28) & (i_3_)) + ((!g1) & (i_5_) & (g28) & (!i_3_)) + ((!g1) & (i_5_) & (g28) & (i_3_)) + ((g1) & (!i_5_) & (!g28) & (!i_3_)) + ((g1) & (!i_5_) & (!g28) & (i_3_)) + ((g1) & (!i_5_) & (g28) & (!i_3_)) + ((g1) & (!i_5_) & (g28) & (i_3_)) + ((g1) & (i_5_) & (!g28) & (!i_3_)) + ((g1) & (i_5_) & (!g28) & (i_3_)) + ((g1) & (i_5_) & (g28) & (!i_3_)) + ((g1) & (i_5_) & (g28) & (i_3_)));
	assign g681 = (((!g1) & (!i_5_) & (!g12) & (i_3_)) + ((!g1) & (i_5_) & (!g12) & (!i_3_)) + ((!g1) & (i_5_) & (!g12) & (i_3_)) + ((!g1) & (i_5_) & (g12) & (!i_3_)) + ((!g1) & (i_5_) & (g12) & (i_3_)) + ((g1) & (!i_5_) & (!g12) & (i_3_)) + ((g1) & (!i_5_) & (g12) & (i_3_)) + ((g1) & (i_5_) & (!g12) & (!i_3_)) + ((g1) & (i_5_) & (!g12) & (i_3_)) + ((g1) & (i_5_) & (g12) & (!i_3_)) + ((g1) & (i_5_) & (g12) & (i_3_)));
	assign g682 = (((!g1) & (!i_5_) & (!g28) & (!i_3_)) + ((!g1) & (!i_5_) & (!g28) & (i_3_)) + ((!g1) & (!i_5_) & (g28) & (!i_3_)) + ((!g1) & (i_5_) & (!g28) & (!i_3_)) + ((!g1) & (i_5_) & (!g28) & (i_3_)) + ((!g1) & (i_5_) & (g28) & (!i_3_)) + ((!g1) & (i_5_) & (g28) & (i_3_)) + ((g1) & (!i_5_) & (!g28) & (!i_3_)) + ((g1) & (!i_5_) & (!g28) & (i_3_)) + ((g1) & (!i_5_) & (g28) & (!i_3_)) + ((g1) & (!i_5_) & (g28) & (i_3_)) + ((g1) & (i_5_) & (!g28) & (!i_3_)) + ((g1) & (i_5_) & (!g28) & (i_3_)) + ((g1) & (i_5_) & (g28) & (!i_3_)) + ((g1) & (i_5_) & (g28) & (i_3_)));
	assign g683 = (((!g684) & (g685)) + ((g684) & (!g685)) + ((g684) & (g685)));
	assign g684 = (((!g27) & (g686)));
	assign g685 = (((g27) & (g689)));
	assign g686 = (((!g687) & (g688)) + ((g687) & (!g688)) + ((g687) & (g688)));
	assign g687 = (((!i_8_) & (g691)));
	assign g688 = (((i_8_) & (g692)));
	assign g689 = (((!i_8_) & (g690)) + ((i_8_) & (!g690)) + ((i_8_) & (g690)));
	assign g690 = (((!i_8_) & (g693)));
	assign g691 = (((!g116) & (!i_7_) & (!g126) & (!i_6_)) + ((!g116) & (!i_7_) & (g126) & (!i_6_)) + ((!g116) & (!i_7_) & (g126) & (i_6_)) + ((!g116) & (i_7_) & (!g126) & (!i_6_)) + ((!g116) & (i_7_) & (!g126) & (i_6_)) + ((!g116) & (i_7_) & (g126) & (!i_6_)) + ((!g116) & (i_7_) & (g126) & (i_6_)) + ((g116) & (!i_7_) & (g126) & (i_6_)) + ((g116) & (i_7_) & (!g126) & (!i_6_)) + ((g116) & (i_7_) & (!g126) & (i_6_)) + ((g116) & (i_7_) & (g126) & (!i_6_)) + ((g116) & (i_7_) & (g126) & (i_6_)));
	assign g692 = (((!g116) & (!i_7_) & (!g5) & (!i_6_)) + ((!g116) & (!i_7_) & (!g5) & (i_6_)) + ((!g116) & (!i_7_) & (g5) & (!i_6_)) + ((!g116) & (!i_7_) & (g5) & (i_6_)) + ((!g116) & (i_7_) & (!g5) & (!i_6_)) + ((!g116) & (i_7_) & (!g5) & (i_6_)) + ((!g116) & (i_7_) & (g5) & (!i_6_)) + ((g116) & (!i_7_) & (!g5) & (i_6_)) + ((g116) & (!i_7_) & (g5) & (i_6_)) + ((g116) & (i_7_) & (!g5) & (!i_6_)) + ((g116) & (i_7_) & (!g5) & (i_6_)) + ((g116) & (i_7_) & (g5) & (!i_6_)));
	assign g693 = (((!i_7_) & (!g126) & (!i_6_)) + ((!i_7_) & (g126) & (!i_6_)) + ((!i_7_) & (g126) & (i_6_)) + ((i_7_) & (!g126) & (!i_6_)) + ((i_7_) & (!g126) & (i_6_)) + ((i_7_) & (g126) & (!i_6_)) + ((i_7_) & (g126) & (i_6_)));
	assign g695 = (((!g47) & (g697)));
	assign g696 = (((g47) & (g699)));
	assign g697 = (((!i_4_) & (g698)) + ((i_4_) & (!g698)) + ((i_4_) & (g698)));
	assign g698 = (((!i_4_) & (g702)));
	assign g699 = (((!g700) & (g701)) + ((g700) & (!g701)) + ((g700) & (g701)));
	assign g700 = (((!i_4_) & (g703)));
	assign g701 = (((i_4_) & (g704)));
	assign g702 = (((!i_5_) & (!g121) & (!i_3_)) + ((!i_5_) & (!g121) & (i_3_)) + ((!i_5_) & (g121) & (!i_3_)) + ((!i_5_) & (g121) & (i_3_)) + ((i_5_) & (!g121) & (!i_3_)) + ((i_5_) & (!g121) & (i_3_)) + ((i_5_) & (g121) & (i_3_)));
	assign g703 = (((!i_5_) & (!g121) & (!i_3_)) + ((!i_5_) & (!g121) & (i_3_)) + ((!i_5_) & (g121) & (!i_3_)) + ((!i_5_) & (g121) & (i_3_)) + ((i_5_) & (!g121) & (!i_3_)) + ((i_5_) & (!g121) & (i_3_)) + ((i_5_) & (g121) & (i_3_)));
	assign g704 = (((!i_6_) & (!i_5_) & (!g27) & (!i_3_)) + ((!i_6_) & (!i_5_) & (g27) & (!i_3_)) + ((!i_6_) & (!i_5_) & (g27) & (i_3_)) + ((!i_6_) & (i_5_) & (!g27) & (!i_3_)) + ((!i_6_) & (i_5_) & (!g27) & (i_3_)) + ((!i_6_) & (i_5_) & (g27) & (!i_3_)) + ((!i_6_) & (i_5_) & (g27) & (i_3_)) + ((i_6_) & (!i_5_) & (!g27) & (!i_3_)) + ((i_6_) & (!i_5_) & (!g27) & (i_3_)) + ((i_6_) & (!i_5_) & (g27) & (!i_3_)) + ((i_6_) & (!i_5_) & (g27) & (i_3_)) + ((i_6_) & (i_5_) & (!g27) & (!i_3_)) + ((i_6_) & (i_5_) & (g27) & (!i_3_)) + ((i_6_) & (i_5_) & (g27) & (i_3_)));
	assign o_1_ = (((!satWreckOut) & (!g82)));
	assign o_2_ = (((!satWreckOut) & (!g199)));
	assign o_3_ = (((!satWreckOut) & (!g263)));
	assign o_4_ = (((!satWreckOut) & (!g320)));
	assign o_5_ = (((!satWreckOut) & (!g356)));
	assign o_6_ = (((!satWreckOut) & (!g395)));
	assign o_7_ = (((!satWreckOut) & (!g418)));
	assign o_8_ = (((!satWreckOut) & (!g437)));
	assign o_9_ = (((!satWreckOut) & (!g454)));
	assign o_10_ = (((!satWreckOut) & (!g467)));
	assign o_11_ = (((!satWreckOut) & (!g490)));
	assign o_12_ = (((!satWreckOut) & (!g510)));
	assign o_13_ = (((!satWreckOut) & (!g520)));
	assign o_14_ = (((!satWreckOut) & (!g523)));
	assign o_15_ = (((!satWreckOut) & (!g532)));
	assign o_16_ = (((!satWreckOut) & (!g537)));
	assign o_17_ = (((!satWreckOut) & (!g540)));
	assign o_18_ = (((!satWreckOut) & (!g542)));
	assign satCompare0 = (((!sk[12]) & (!sk[13]) & (!sk[14]) & (!i_0_) & (!i_1_) & (!i_2_)) + ((!sk[12]) & (!sk[13]) & (sk[14]) & (!i_0_) & (!i_1_) & (i_2_)) + ((!sk[12]) & (sk[13]) & (!sk[14]) & (!i_0_) & (i_1_) & (!i_2_)) + ((!sk[12]) & (sk[13]) & (sk[14]) & (!i_0_) & (i_1_) & (i_2_)) + ((sk[12]) & (!sk[13]) & (!sk[14]) & (i_0_) & (!i_1_) & (!i_2_)) + ((sk[12]) & (!sk[13]) & (sk[14]) & (i_0_) & (!i_1_) & (i_2_)) + ((sk[12]) & (sk[13]) & (!sk[14]) & (i_0_) & (i_1_) & (!i_2_)) + ((sk[12]) & (sk[13]) & (sk[14]) & (i_0_) & (i_1_) & (i_2_)));
	assign satCompare1 = (((!sk[15]) & (!sk[16]) & (!sk[17]) & (!i_6_) & (!i_7_) & (!i_8_)) + ((!sk[15]) & (!sk[16]) & (sk[17]) & (!i_6_) & (!i_7_) & (i_8_)) + ((!sk[15]) & (sk[16]) & (!sk[17]) & (!i_6_) & (i_7_) & (!i_8_)) + ((!sk[15]) & (sk[16]) & (sk[17]) & (!i_6_) & (i_7_) & (i_8_)) + ((sk[15]) & (!sk[16]) & (!sk[17]) & (i_6_) & (!i_7_) & (!i_8_)) + ((sk[15]) & (!sk[16]) & (sk[17]) & (i_6_) & (!i_7_) & (i_8_)) + ((sk[15]) & (sk[16]) & (!sk[17]) & (i_6_) & (i_7_) & (!i_8_)) + ((sk[15]) & (sk[16]) & (sk[17]) & (i_6_) & (i_7_) & (i_8_)));
	assign satCompare2 = (((!sk[18]) & (!sk[19]) & (!sk[20]) & (!i_3_) & (!i_4_) & (!i_5_)) + ((!sk[18]) & (!sk[19]) & (sk[20]) & (!i_3_) & (!i_4_) & (i_5_)) + ((!sk[18]) & (sk[19]) & (!sk[20]) & (!i_3_) & (i_4_) & (!i_5_)) + ((!sk[18]) & (sk[19]) & (sk[20]) & (!i_3_) & (i_4_) & (i_5_)) + ((sk[18]) & (!sk[19]) & (!sk[20]) & (i_3_) & (!i_4_) & (!i_5_)) + ((sk[18]) & (!sk[19]) & (sk[20]) & (i_3_) & (!i_4_) & (i_5_)) + ((sk[18]) & (sk[19]) & (!sk[20]) & (i_3_) & (i_4_) & (!i_5_)) + ((sk[18]) & (sk[19]) & (sk[20]) & (i_3_) & (i_4_) & (i_5_)));
	assign satCompareLevel0_0 = (((satCompare0) & (satCompare1) & (satCompare2)));
	assign satMask0 = (((!sk[12]) & (!sk[13]) & (sk[14]) & (sk[15]) & (sk[16]) & (sk[17])));
	assign satMask1 = (((sk[18]) & (!sk[19]) & (sk[20])));
	assign satMaskLevel0_0 = (((satMask0) & (satMask1)));
	assign satWreckOut = (((satCompareLevel0_0) & (!satMaskLevel0_0)));
endmodule
