module seqx6xv (i_40_, i_30_, i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_, i_4_, i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_, i_16_, i_22_, i_15_, i_32_, i_31_, i_34_, i_33_, i_19_, i_36_, i_35_, i_38_, i_29_, i_37_, o_1_, o_19_, o_2_, o_0_, o_29_, o_25_, o_12_, o_26_, o_11_, o_27_, o_14_, o_28_, o_13_, o_34_, o_21_, o_16_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_, o_31_, o_24_, o_17_, o_30_, o_20_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

	input i_40_;
	input i_30_;
	input i_20_;
	input i_9_;
	input i_10_;
	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_27_;
	input i_14_;
	input i_3_;
	input i_39_;
	input i_28_;
	input i_13_;
	input i_4_;
	input i_25_;
	input i_12_;
	input i_1_;
	input i_26_;
	input i_11_;
	input i_2_;
	input i_23_;
	input i_18_;
	input i_24_;
	input i_17_;
	input i_0_;
	input i_21_;
	input i_16_;
	input i_22_;
	input i_15_;
	input i_32_;
	input i_31_;
	input i_34_;
	input i_33_;
	input i_19_;
	input i_36_;
	input i_35_;
	input i_38_;
	input i_29_;
	input i_37_;
	output o_1_;
	output o_19_;
	output o_2_;
	output o_0_;
	output o_29_;
	output o_25_;
	output o_12_;
	output o_26_;
	output o_11_;
	output o_27_;
	output o_14_;
	output o_28_;
	output o_13_;
	output o_34_;
	output o_21_;
	output o_16_;
	output o_33_;
	output o_22_;
	output o_15_;
	output o_32_;
	output o_23_;
	output o_18_;
	output o_31_;
	output o_24_;
	output o_17_;
	output o_30_;
	output o_20_;
	output o_10_;
	output o_9_;
	output o_7_;
	output o_8_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;

	wire [1064 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], x6758x, n_n1135, n_n1134, x6747x, x6757x}, o_1_);
	defparam lut_3.LUT_SIZE = 6;
	defparam lut_3.mask = 64'h3f3fffff7fffffff;

	lut_sub lut_9 ({sk[1], i_6_, i_36_, x6771x, x1874x, x313x, n_n866}, o_19_);
	defparam lut_9.LUT_SIZE = 7;
	defparam lut_9.mask = 128'h5f5f5f5f5f5f5f5f00ff00ff0fff1fff;

	lut_sub lut_13 ({sk[2], n_n1165, x6806x, x6807x, x6808x}, o_2_);
	defparam lut_13.LUT_SIZE = 5;
	defparam lut_13.mask = 32'h5f5f7fff;

	lut_sub lut_18 ({sk[3], x6929x, x6916x, n_n1094, n_n1088, n_n1086, x6904x}, o_0_);
	defparam lut_18.LUT_SIZE = 7;
	defparam lut_18.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_25 ({sk[4], x6937x, x366x, x529x, n_n1935, n_n1965, n_n1993}, o_29_);
	defparam lut_25.LUT_SIZE = 7;
	defparam lut_25.mask = 128'h77777f7f77777f7f7f7f7fffffffffff;

	lut_sub lut_31 ({sk[5], n_n1581, x6965x, x6966x, x6982x, x6983x, x6987x}, o_25_);
	defparam lut_31.LUT_SIZE = 7;
	defparam lut_31.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_38 ({sk[6], i_40_, i_7_, i_8_, i_5_, i_0_, x554x}, o_12_);
	defparam lut_38.LUT_SIZE = 7;
	defparam lut_38.mask = 128'h77777f7f77777f7f0004000000000000;

	lut_sub lut_40 ({sk[7], x7005x, x6998x, x238x, x6994x}, o_26_);
	defparam lut_40.LUT_SIZE = 5;
	defparam lut_40.mask = 32'h00ff7fff;

	lut_sub lut_45 ({sk[8], x7023x, n_n1014, x1626x, n_n1009, x1630x, x7012x}, o_11_);
	defparam lut_45.LUT_SIZE = 7;
	defparam lut_45.mask = 128'h77777f7f77777f7f00ff07ffffffffff;

	lut_sub lut_50 ({sk[9], x6982x, x6983x, n_n1628, n_n1630, n_n1631, x7038x}, o_27_);
	defparam lut_50.LUT_SIZE = 7;
	defparam lut_50.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_57 ({sk[10], i_13_, o_15_, n_n973, x51x, n_n967, x530x}, o_14_);
	defparam lut_57.LUT_SIZE = 7;
	defparam lut_57.mask = 128'h77777f7f77777f7f030fffff575fffff;

	lut_sub lut_62 ({sk[11], n_n1011, x335x, x373x, x396x, n_n1971, x89x}, o_28_);
	defparam lut_62.LUT_SIZE = 7;
	defparam lut_62.mask = 128'h77777f7f77777f7f33373f3f37373f3f;

	lut_sub lut_67 ({sk[12], i_40_, i_39_, i_38_, o_15_, x391x, x51x}, o_13_);
	defparam lut_67.LUT_SIZE = 7;
	defparam lut_67.mask = 128'h77777f7f77777f7f3f5f0f0f3f0f5f0f;

	lut_sub lut_72 ({sk[13], n_n1716, x7072x, n_n1715, x7093x, x7094x}, o_34_);
	defparam lut_72.LUT_SIZE = 6;
	defparam lut_72.mask = 64'h55ffffff7fffffff;

	lut_sub lut_78 ({sk[14], x1518x, x1519x, x1505x, x1506x, x7110x}, o_21_);
	defparam lut_78.LUT_SIZE = 6;
	defparam lut_78.mask = 64'h55ffffff7fffffff;

	lut_sub lut_84 ({sk[15], x411x, x436x, x1498x, x7117x, x7118x}, o_16_);
	defparam lut_84.LUT_SIZE = 6;
	defparam lut_84.mask = 64'h55ffffff7f7f7fff;

	lut_sub lut_89 ({sk[16], x7140x, x7141x, x7185x, x7186x, x8533x}, o_33_);
	defparam lut_89.LUT_SIZE = 6;
	defparam lut_89.mask = 64'h55ffffffbfffffff;

	lut_sub lut_95 ({sk[17], n_n967, x1391x, n_n1531, n_n673, x7203x, x7223x}, o_22_);
	defparam lut_95.LUT_SIZE = 7;
	defparam lut_95.mask = 128'h77777f7f77777f7f77ffffff7fffffff;

	lut_sub lut_101 ({sk[18], i_7_, i_33_}, o_15_);
	defparam lut_101.LUT_SIZE = 3;
	defparam lut_101.mask = 8'h31;

	lut_sub lut_103 ({sk[19], i_40_, i_7_, i_32_, i_33_, n_n979, n_n1005}, o_32_);
	defparam lut_103.LUT_SIZE = 7;
	defparam lut_103.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_105 ({sk[20], x7272x, x7251x, x7249x, x7250x, x7269x, x7270x}, o_23_);
	defparam lut_105.LUT_SIZE = 7;
	defparam lut_105.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_112 ({sk[21], x7346x, x7301x, x7302x}, o_18_);
	defparam lut_112.LUT_SIZE = 4;
	defparam lut_112.mask = 16'h157f;

	lut_sub lut_116 ({sk[22], n_n837, x54x, n_n1908, n_n1907, x7358x, x8563x}, o_31_);
	defparam lut_116.LUT_SIZE = 7;
	defparam lut_116.mask = 128'h77777f7f77777f7fbfffbfffbfffffff;

	lut_sub lut_122 ({sk[23], n_n2581, x6982x, x6983x, n_n2838, x7386x, x7383x}, o_24_);
	defparam lut_122.LUT_SIZE = 7;
	defparam lut_122.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_129 ({sk[24], n_n1409, n_n1414, n_n1412, x7412x, x7448x}, o_17_);
	defparam lut_129.LUT_SIZE = 6;
	defparam lut_129.mask = 64'h55ffffff7fffffff;

	lut_sub lut_135 ({sk[25], i_24_, x415x, x423x, n_n1651, x7463x}, o_30_);
	defparam lut_135.LUT_SIZE = 6;
	defparam lut_135.mask = 64'h55ffffff77777fff;

	lut_sub lut_140 ({sk[26], n_n1484, x7494x, x7495x, n_n1489, x7506x}, o_20_);
	defparam lut_140.LUT_SIZE = 6;
	defparam lut_140.mask = 64'h55ffffff7fffffff;

	lut_sub lut_146 ({sk[27], n_n1384, n_n982, x328x, x325x, x1031x, x1032x}, o_10_);
	defparam lut_146.LUT_SIZE = 7;
	defparam lut_146.mask = 128'h77777f7f77777f7f777f77ffffffffff;

	lut_sub lut_152 ({sk[28], x7530x, x109x, n_n1372, n_n1048, n_n785, x7526x}, o_9_);
	defparam lut_152.LUT_SIZE = 7;
	defparam lut_152.mask = 128'h77777f7f77777f7f55ff57ffffffffff;

	lut_sub lut_157 ({sk[29], n_n1375, n_n1374, n_n1356, x7546x, x7547x}, o_7_);
	defparam lut_157.LUT_SIZE = 6;
	defparam lut_157.mask = 64'h55ffffff7fffffff;

	lut_sub lut_163 ({sk[30], i_7_, i_33_, i_38_, n_n1064, x146x, x340x}, o_8_);
	defparam lut_163.LUT_SIZE = 7;
	defparam lut_163.mask = 128'h77777f7f77777f7f333733373337ffff;

	lut_sub lut_167 ({sk[31], x7639x, x7616x, n_n1280, n_n1282, x7574x, x7615x}, o_5_);
	defparam lut_167.LUT_SIZE = 7;
	defparam lut_167.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_174 ({sk[32], x7684x, x536x, n_n1329, x7674x}, o_6_);
	defparam lut_174.LUT_SIZE = 5;
	defparam lut_174.mask = 32'h00ff7fff;

	lut_sub lut_179 ({sk[33], x7732x, n_n1184, n_n1197, x7730x, x7763x, x7764x}, o_3_);
	defparam lut_179.LUT_SIZE = 7;
	defparam lut_179.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_186 ({sk[34], x7824x, n_n785, x483x, x7820x, x463x, x7821x}, o_4_);
	defparam lut_186.LUT_SIZE = 7;
	defparam lut_186.mask = 128'h77777f7f77777f7f55557fffffffffff;

	lut_sub lut_192 ({sk[35], x1923x, x6726x, x145x, x1883x, x6752x}, x6758x);
	defparam lut_192.LUT_SIZE = 6;
	defparam lut_192.mask = 64'h55ffffff7fffffff;

	lut_sub lut_198 ({sk[36], i_32_, x525x, x347x, x1913x, x1912x, x6733x}, n_n1135);
	defparam lut_198.LUT_SIZE = 7;
	defparam lut_198.mask = 128'h77777f7f77777f7f7f7f7fff7f7f7f7f;

	lut_sub lut_203 ({sk[37], i_5_, i_37_, n_n1011, x353x, x6740x, x6741x}, n_n1134);
	defparam lut_203.LUT_SIZE = 7;
	defparam lut_203.mask = 128'h77777f7f77777f7f7f7f7f7777777777;

	lut_sub lut_208 ({sk[38], n_n1074, n_n560, n_n884, x303x, x6745x, x6746x}, x6747x);
	defparam lut_208.LUT_SIZE = 7;
	defparam lut_208.mask = 128'h77777f7f77777f7f557f557f557f55ff;

	lut_sub lut_213 ({sk[39], x1934x, n_n1001, n_n975, n_n905, x6718x, x8546x}, x6757x);
	defparam lut_213.LUT_SIZE = 7;
	defparam lut_213.mask = 128'h77777f7f77777f7fbbbfbfbfffffffff;

	lut_sub lut_219 ({sk[40], n_n985, n_n515, n_n1008, x1867x, x6767x, x6768x}, x6771x);
	defparam lut_219.LUT_SIZE = 7;
	defparam lut_219.mask = 128'h77777f7f77777f7f7f7f7f7f7f7f7fff;

	lut_sub lut_224 ({sk[41], i_7_, n_n1014, n_n1061, x50x, x80x, n_n582}, x1874x);
	defparam lut_224.LUT_SIZE = 7;
	defparam lut_224.mask = 128'h77777f7f77777f7f0000111f00000000;

	lut_sub lut_227 ({sk[42], i_7_, i_32_, i_34_, i_33_, i_35_}, x313x);
	defparam lut_227.LUT_SIZE = 6;
	defparam lut_227.mask = 64'h55ffffff10000000;

	lut_sub lut_229 ({sk[43], i_40_, i_38_, i_37_}, n_n866);
	defparam lut_229.LUT_SIZE = 4;
	defparam lut_229.mask = 16'h1504;

	lut_sub lut_231 ({sk[44], x1844x, x1846x, x6793x, x6794x}, n_n1165);
	defparam lut_231.LUT_SIZE = 5;
	defparam lut_231.mask = 32'h00ff7fff;

	lut_sub lut_236 ({sk[45], i_10_, n_n982, n_n1164, x397x, x8545x, x8551x}, x6806x);
	defparam lut_236.LUT_SIZE = 7;
	defparam lut_236.mask = 128'h77777f7f77777f7feeffefffeeffeeff;

	lut_sub lut_241 ({sk[46], x145x, n_n1373, x72x, x432x, x491x, x6803x}, x6807x);
	defparam lut_241.LUT_SIZE = 7;
	defparam lut_241.mask = 128'h77777f7f77777f7f5557ffffffffffff;

	lut_sub lut_246 ({sk[47], x48x, x247x, x1831x, x52x, n_n1072, x42x}, x6808x);
	defparam lut_246.LUT_SIZE = 7;
	defparam lut_246.mask = 128'h77777f7f77777f7f0000ffff01ffffff;

	lut_sub lut_250 ({sk[48], n_n1083, n_n1084, x1706x, x6922x, x6923x, x8544x}, x6929x);
	defparam lut_250.LUT_SIZE = 7;
	defparam lut_250.mask = 128'h77777f7f77777f7fbfffffffffffffff;

	lut_sub lut_257 ({sk[49], n_n1093, n_n1091, x6879x, x6878x, x6913x}, x6916x);
	defparam lut_257.LUT_SIZE = 6;
	defparam lut_257.mask = 64'h55ffffff7fffffff;

	lut_sub lut_263 ({sk[50], i_23_, x1791x, x1792x, x1789x}, n_n1094);
	defparam lut_263.LUT_SIZE = 5;
	defparam lut_263.mask = 32'h00ff7f55;

	lut_sub lut_267 ({sk[51], i_24_, x50x, x54x, x87x, x1751x, x8562x}, n_n1088);
	defparam lut_267.LUT_SIZE = 7;
	defparam lut_267.mask = 128'h77777f7f77777f7fbbbbbbbfbbbbbbbb;

	lut_sub lut_271 ({sk[52], x431x, x541x, x227x, x149x, x155x, x6892x}, n_n1086);
	defparam lut_271.LUT_SIZE = 7;
	defparam lut_271.mask = 128'h77777f7f77777f7f7fff7fff7fffffff;

	lut_sub lut_277 ({sk[53], x541x, x362x, x148x, n_n1108, x1731x, x6901x}, x6904x);
	defparam lut_277.LUT_SIZE = 7;
	defparam lut_277.mask = 128'h77777f7f77777f7f7fff7fff7fffffff;

	lut_sub lut_283 ({sk[54], i_21_, i_15_, x35x, n_n1936, x552x, x1694x}, x6937x);
	defparam lut_283.LUT_SIZE = 7;
	defparam lut_283.mask = 128'h77777f7f77777f7f5f5f5f7f5f5f5f5f;

	lut_sub lut_287 ({sk[55], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x366x);
	defparam lut_287.LUT_SIZE = 7;
	defparam lut_287.mask = 128'h77777f7f77777f7f0000400000000000;

	lut_sub lut_289 ({sk[56], i_32_, i_31_, i_34_, i_33_, x6834x}, x529x);
	defparam lut_289.LUT_SIZE = 6;
	defparam lut_289.mask = 64'h55ffffff10000000;

	lut_sub lut_291 ({sk[57], i_40_, i_39_, i_36_, i_35_, i_38_, x529x}, n_n1935);
	defparam lut_291.LUT_SIZE = 7;
	defparam lut_291.mask = 128'h77777f7f77777f7f0000000010000000;

	lut_sub lut_293 ({sk[58], i_31_, i_37_, n_n1074, n_n964, n_n799, x6862x}, n_n1965);
	defparam lut_293.LUT_SIZE = 7;
	defparam lut_293.mask = 128'h77777f7f77777f7f0000000100000000;

	lut_sub lut_295 ({sk[59], i_40_, i_7_, i_32_, i_33_, n_n1002, n_n795}, n_n1993);
	defparam lut_295.LUT_SIZE = 7;
	defparam lut_295.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_297 ({sk[60], x1691x, x1692x, x6940x, x6941x, x6942x}, n_n1581);
	defparam lut_297.LUT_SIZE = 6;
	defparam lut_297.mask = 64'h55ffffff7fffffff;

	lut_sub lut_303 ({sk[61], x1682x, x6946x, n_n1118, x1675x, x6950x, x6951x}, x6965x);
	defparam lut_303.LUT_SIZE = 7;
	defparam lut_303.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_310 ({sk[62], n_n833, n_n764, x240x, n_n1908, n_n1907, x8542x}, x6966x);
	defparam lut_310.LUT_SIZE = 7;
	defparam lut_310.mask = 128'h77777f7f77777f7fbfffbfffbfffffff;

	lut_sub lut_316 ({sk[63], x82x, n_n1048, n_n785, x87x, x37x, x1653x}, x6982x);
	defparam lut_316.LUT_SIZE = 7;
	defparam lut_316.mask = 128'h77777f7f77777f7f5555555d555555dd;

	lut_sub lut_320 ({sk[64], x1652x, x1661x, x6970x, x6971x, x8541x}, x6983x);
	defparam lut_320.LUT_SIZE = 6;
	defparam lut_320.mask = 64'h55ffffffbfffffff;

	lut_sub lut_326 ({sk[65], x335x, n_n2581, x396x, n_n1971, x173x, x181x}, x6987x);
	defparam lut_326.LUT_SIZE = 7;
	defparam lut_326.mask = 128'h77777f7f77777f7f7f7fffff7fffffff;

	lut_sub lut_332 ({sk[66], i_34_, i_36_, i_35_, i_38_, i_37_, x46x}, x554x);
	defparam lut_332.LUT_SIZE = 7;
	defparam lut_332.mask = 128'h77777f7f77777f7f0000000140000000;

	lut_sub lut_335 ({sk[67], x429x, n_n2838, n_n2836, x71x, x302x, x8540x}, x7005x);
	defparam lut_335.LUT_SIZE = 7;
	defparam lut_335.mask = 128'h77777f7f77777f7fabffffffafffffff;

	lut_sub lut_341 ({sk[68], i_3_, i_4_, i_1_, x314x, n_n926, n_n833}, x6998x);
	defparam lut_341.LUT_SIZE = 7;
	defparam lut_341.mask = 128'h77777f7f77777f7f0005050507070707;

	lut_sub lut_346 ({sk[69], i_7_, i_39_, i_2_, n_n985, n_n833, x80x}, x238x);
	defparam lut_346.LUT_SIZE = 7;
	defparam lut_346.mask = 128'h77777f7f77777f7f0015001100000000;

	lut_sub lut_349 ({sk[70], i_4_, i_1_, i_0_, x431x, x436x, x79x}, x6994x);
	defparam lut_349.LUT_SIZE = 7;
	defparam lut_349.mask = 128'h77777f7f77777f7f0011001100150005;

	lut_sub lut_353 ({sk[71], n_n926, x92x, x319x, x470x, x7018x, x7021x}, x7023x);
	defparam lut_353.LUT_SIZE = 7;
	defparam lut_353.mask = 128'h77777f7f77777f7f5555555f777f777f;

	lut_sub lut_358 ({sk[72], i_40_, i_39_}, n_n1014);
	defparam lut_358.LUT_SIZE = 3;
	defparam lut_358.mask = 8'h31;

	lut_sub lut_360 ({sk[73], i_9_, i_12_, i_11_, x47x, x341x, x412x}, x1626x);
	defparam lut_360.LUT_SIZE = 7;
	defparam lut_360.mask = 128'h77777f7f77777f7f1111111111131313;

	lut_sub lut_364 ({sk[74], i_36_, i_38_, i_37_}, n_n1009);
	defparam lut_364.LUT_SIZE = 4;
	defparam lut_364.mask = 16'h1520;

	lut_sub lut_366 ({sk[75], i_15_, n_n1066, n_n860, n_n933, x39x, x1633x}, x1630x);
	defparam lut_366.LUT_SIZE = 7;
	defparam lut_366.mask = 128'h77777f7f77777f7f0000005500000057;

	lut_sub lut_369 ({sk[76], i_9_, i_11_, x47x, x319x, x78x, x388x}, x7012x);
	defparam lut_369.LUT_SIZE = 7;
	defparam lut_369.mask = 128'h77777f7f77777f7f0003000000130000;

	lut_sub lut_372 ({sk[77], i_40_, x173x, x181x, n_n837, n_n836, x6946x}, n_n1628);
	defparam lut_372.LUT_SIZE = 7;
	defparam lut_372.mask = 128'h77777f7f77777f7f55ffffff57ffffff;

	lut_sub lut_377 ({sk[78], x7028x, n_n1980, x68x, x504x, x157x}, n_n1630);
	defparam lut_377.LUT_SIZE = 6;
	defparam lut_377.mask = 64'h55ffffff57ffffff;

	lut_sub lut_382 ({sk[79], n_n1927, n_n2793, n_n2456, x300x, x8539x}, n_n1631);
	defparam lut_382.LUT_SIZE = 6;
	defparam lut_382.mask = 64'h55ffffffbfffffff;

	lut_sub lut_388 ({sk[80], n_n1928, n_n1983, n_n837, x54x, x7034x, x8558x}, x7038x);
	defparam lut_388.LUT_SIZE = 7;
	defparam lut_388.mask = 128'h77777f7f77777f7fbbbfffffffffffff;

	lut_sub lut_394 ({sk[81], i_40_, i_39_, i_38_}, n_n973);
	defparam lut_394.LUT_SIZE = 4;
	defparam lut_394.mask = 16'h1502;

	lut_sub lut_396 ({sk[82], i_32_, i_34_, i_33_, i_36_, i_35_, i_37_}, x51x);
	defparam lut_396.LUT_SIZE = 7;
	defparam lut_396.mask = 128'h77777f7f77777f7f0020000000000000;

	lut_sub lut_398 ({sk[83], i_40_, i_39_, i_38_}, n_n967);
	defparam lut_398.LUT_SIZE = 4;
	defparam lut_398.mask = 16'h1540;

	lut_sub lut_400 ({sk[84], i_39_, i_32_, i_33_, i_38_, i_37_, n_n1002}, x530x);
	defparam lut_400.LUT_SIZE = 7;
	defparam lut_400.mask = 128'h77777f7f77777f7f0040000000000000;

	lut_sub lut_402 ({sk[85], i_39_, i_38_}, n_n1011);
	defparam lut_402.LUT_SIZE = 3;
	defparam lut_402.mask = 8'h38;

	lut_sub lut_404 ({sk[86], i_36_, i_35_, i_38_, i_37_, n_n1074}, x335x);
	defparam lut_404.LUT_SIZE = 6;
	defparam lut_404.mask = 64'h55ffffff00000001;

	lut_sub lut_406 ({sk[87], i_40_, i_38_}, x373x);
	defparam lut_406.LUT_SIZE = 3;
	defparam lut_406.mask = 8'h38;

	lut_sub lut_408 ({sk[88], i_7_, i_3_, i_4_, i_1_, i_2_, i_0_}, x396x);
	defparam lut_408.LUT_SIZE = 7;
	defparam lut_408.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_410 ({sk[89], i_40_, i_7_, i_39_, i_38_, n_n1074, x6895x}, n_n1971);
	defparam lut_410.LUT_SIZE = 7;
	defparam lut_410.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_412 ({sk[90], i_32_, i_34_, i_33_, i_36_, i_35_, i_37_}, x89x);
	defparam lut_412.LUT_SIZE = 7;
	defparam lut_412.mask = 128'h77777f7f77777f7f0000008000000000;

	lut_sub lut_414 ({sk[91], i_32_, i_34_, i_33_, i_36_, i_35_, i_37_}, x391x);
	defparam lut_414.LUT_SIZE = 7;
	defparam lut_414.mask = 128'h77777f7f77777f7f0002000000000000;

	lut_sub lut_416 ({sk[92], i_1_, i_2_, i_0_, x518x, x1567x, x7061x}, n_n1716);
	defparam lut_416.LUT_SIZE = 7;
	defparam lut_416.mask = 128'h77777f7f77777f7f777f777777777777;

	lut_sub lut_420 ({sk[93], x1575x, x1557x, x7069x, x8538x}, x7072x);
	defparam lut_420.LUT_SIZE = 5;
	defparam lut_420.mask = 32'h00ffbfff;

	lut_sub lut_425 ({sk[94], x387x, x119x, x1538x, x7084x, x7085x}, n_n1715);
	defparam lut_425.LUT_SIZE = 6;
	defparam lut_425.mask = 64'h55ffffff7f7f7fff;

	lut_sub lut_430 ({sk[95], i_37_, n_n1011, x7048x, x424x, x1583x, x7092x}, x7093x);
	defparam lut_430.LUT_SIZE = 7;
	defparam lut_430.mask = 128'h77777f7f77777f7f7fff7fff7fff77ff;

	lut_sub lut_436 ({sk[96], n_n1074, x817x, x1524x, x7075x, x7076x}, x7094x);
	defparam lut_436.LUT_SIZE = 6;
	defparam lut_436.mask = 64'h55ffffff7f7f7fff;

	lut_sub lut_441 ({sk[97], i_7_, i_6_, i_34_, i_38_, n_n1014, n_n864}, x1518x);
	defparam lut_441.LUT_SIZE = 7;
	defparam lut_441.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_443 ({sk[98], i_0_, n_n991, x47x, x453x, x436x, x400x}, x1519x);
	defparam lut_443.LUT_SIZE = 7;
	defparam lut_443.mask = 128'h77777f7f77777f7f0303035700000000;

	lut_sub lut_446 ({sk[99], i_0_, n_n1002, x47x, x7104x, x100x, x1514x}, x1505x);
	defparam lut_446.LUT_SIZE = 7;
	defparam lut_446.mask = 128'h77777f7f77777f7f005f007f00000000;

	lut_sub lut_450 ({sk[100], i_7_, i_6_, i_34_, x1510x, n_n1072, n_n1012}, x1506x);
	defparam lut_450.LUT_SIZE = 7;
	defparam lut_450.mask = 128'h77777f7f77777f7f0f1f0f0f00000000;

	lut_sub lut_453 ({sk[101], i_6_, i_33_, i_35_, n_n978, x355x, x453x}, x7110x);
	defparam lut_453.LUT_SIZE = 7;
	defparam lut_453.mask = 128'h77777f7f77777f7fffff0001ffff0000;

	lut_sub lut_456 ({sk[102], i_1_, i_2_, i_0_, n_n1074, n_n842}, x411x);
	defparam lut_456.LUT_SIZE = 6;
	defparam lut_456.mask = 64'h55ffffff00000100;

	lut_sub lut_458 ({sk[103], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x436x);
	defparam lut_458.LUT_SIZE = 7;
	defparam lut_458.mask = 128'h77777f7f77777f7f0004000000000000;

	lut_sub lut_460 ({sk[104], i_39_, i_38_, i_37_, x88x, n_n991, x528x}, x1498x);
	defparam lut_460.LUT_SIZE = 7;
	defparam lut_460.mask = 128'h77777f7f77777f7f0000005700000000;

	lut_sub lut_463 ({sk[105], n_n861, n_n991, n_n880, n_n975, n_n971, x390x}, x7117x);
	defparam lut_463.LUT_SIZE = 7;
	defparam lut_463.mask = 128'h77777f7f77777f7f0011001100110f1f;

	lut_sub lut_466 ({sk[106], n_n970, x362x, n_n997, x510x, x526x, x346x}, x7118x);
	defparam lut_466.LUT_SIZE = 7;
	defparam lut_466.mask = 128'h77777f7f77777f7f000f333f111f333f;

	lut_sub lut_470 ({sk[107], x52x, n_n1375, x7134x, x36x, x1476x, x7135x}, x7140x);
	defparam lut_470.LUT_SIZE = 7;
	defparam lut_470.mask = 128'h77777f7f77777f7f7777ffff777fffff;

	lut_sub lut_475 ({sk[108], n_n937, n_n1374, x386x, x1489x, x7129x, x1475x}, x7141x);
	defparam lut_475.LUT_SIZE = 7;
	defparam lut_475.mask = 128'h77777f7f77777f7f7f7fffff7fffffff;

	lut_sub lut_481 ({sk[109], x342x, n_n905, x1467x, x1466x, x7143x, x7183x}, x7185x);
	defparam lut_481.LUT_SIZE = 7;
	defparam lut_481.mask = 128'h77777f7f77777f7f7fff7fff7fffffff;

	lut_sub lut_487 ({sk[110], i_36_, n_n960, x7152x, x812x, x1460x, x1461x}, x7186x);
	defparam lut_487.LUT_SIZE = 7;
	defparam lut_487.mask = 128'h77777f7f77777f7f77ff7fff77ff77ff;

	lut_sub lut_492 ({sk[111], i_32_, i_33_, x122x, n_n1675, x7176x, x7175x}, x8533x);
	defparam lut_492.LUT_SIZE = 7;
	defparam lut_492.mask = 128'h77777f7f77777f7f8000800000008000;

	lut_sub lut_495 ({sk[112], i_31_, i_38_, i_37_, x49x, n_n673, x8571x}, x1391x);
	defparam lut_495.LUT_SIZE = 7;
	defparam lut_495.mask = 128'h77777f7f77777f7f3b00000033000000;

	lut_sub lut_498 ({sk[113], n_n973, x362x, x7210x, x428x, n_n673, x1383x}, n_n1531);
	defparam lut_498.LUT_SIZE = 7;
	defparam lut_498.mask = 128'h77777f7f77777f7f55ff5fff77ff7fff;

	lut_sub lut_503 ({sk[114], i_12_, i_16_, i_15_, i_31_, x49x}, n_n673);
	defparam lut_503.LUT_SIZE = 6;
	defparam lut_503.mask = 64'h55ffffff00000004;

	lut_sub lut_505 ({sk[115], i_35_, i_37_, n_n883, n_n977, x301x, x428x}, x7203x);
	defparam lut_505.LUT_SIZE = 7;
	defparam lut_505.mask = 128'h77777f7f77777f7f3333337733333737;

	lut_sub lut_509 ({sk[116], i_14_, i_15_, x405x, x41x, x7222x, x8532x}, x7223x);
	defparam lut_509.LUT_SIZE = 7;
	defparam lut_509.mask = 128'h77777f7f77777f7fbbffbbffbbffbbbf;

	lut_sub lut_515 ({sk[117], i_34_, i_36_, i_35_}, n_n979);
	defparam lut_515.LUT_SIZE = 4;
	defparam lut_515.mask = 16'h1540;

	lut_sub lut_517 ({sk[118], i_39_, i_38_, i_37_}, n_n1005);
	defparam lut_517.LUT_SIZE = 4;
	defparam lut_517.mask = 16'h1510;

	lut_sub lut_519 ({sk[119], x7237x, x7261x, x1356x, x7260x, x8531x}, x7272x);
	defparam lut_519.LUT_SIZE = 6;
	defparam lut_519.mask = 64'h55ffffffbfffffff;

	lut_sub lut_525 ({sk[120], i_40_, i_39_, i_35_, i_38_, i_37_, n_n1074}, x7251x);
	defparam lut_525.LUT_SIZE = 7;
	defparam lut_525.mask = 128'h77777f7f77777f7f0000001400000000;

	lut_sub lut_528 ({sk[121], i_0_, i_32_, i_33_, x373x, n_n715, x336x}, x7249x);
	defparam lut_528.LUT_SIZE = 7;
	defparam lut_528.mask = 128'h77777f7f77777f7f5555555555575555;

	lut_sub lut_531 ({sk[122], i_40_, i_39_, i_38_, n_n966, n_n1012, x1341x}, x7250x);
	defparam lut_531.LUT_SIZE = 7;
	defparam lut_531.mask = 128'h77777f7f77777f7f5555575557555755;

	lut_sub lut_535 ({sk[123], i_40_, n_n1009, n_n874, n_n462, x7266x, x7267x}, x7269x);
	defparam lut_535.LUT_SIZE = 7;
	defparam lut_535.mask = 128'h77777f7f77777f7f777f777f777f77ff;

	lut_sub lut_540 ({sk[124], x1364x, x1349x, x7243x, x7244x, x8530x}, x7270x);
	defparam lut_540.LUT_SIZE = 6;
	defparam lut_540.mask = 64'h55ffffffbfffffff;

	lut_sub lut_546 ({sk[125], x7329x, n_n1447, n_n1453, n_n1452, x7344x}, x7346x);
	defparam lut_546.LUT_SIZE = 6;
	defparam lut_546.mask = 64'h55ffffff7fffffff;

	lut_sub lut_552 ({sk[126], x1308x, x7283x, x7284x, x7299x, x8526x}, x7301x);
	defparam lut_552.LUT_SIZE = 6;
	defparam lut_552.mask = 64'h55ffffffbfffffff;

	lut_sub lut_558 ({sk[127], i_40_, x764x, x1284x, x1285x, x1293x, x1294x}, x7302x);
	defparam lut_558.LUT_SIZE = 7;
	defparam lut_558.mask = 128'h77777f7f77777f7f7fffffff7fff7fff;

	lut_sub lut_564 ({sk[128], i_24_, i_32_, i_34_, i_33_, i_35_, x82x}, n_n837);
	defparam lut_564.LUT_SIZE = 7;
	defparam lut_564.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_566 ({sk[129], i_39_, i_36_, i_38_, i_37_}, x54x);
	defparam lut_566.LUT_SIZE = 5;
	defparam lut_566.mask = 32'h00ff8020;

	lut_sub lut_569 ({sk[130], i_40_, i_38_, n_n842, x89x, n_n843}, n_n1908);
	defparam lut_569.LUT_SIZE = 6;
	defparam lut_569.mask = 64'h55ffffff01000000;

	lut_sub lut_571 ({sk[131], i_39_, i_38_, n_n842, x89x, n_n843}, n_n1907);
	defparam lut_571.LUT_SIZE = 6;
	defparam lut_571.mask = 64'h55ffffff01000000;

	lut_sub lut_573 ({sk[132], i_40_, n_n1971, n_n837, x245x, n_n836, x8565x}, x7358x);
	defparam lut_573.LUT_SIZE = 7;
	defparam lut_573.mask = 128'h77777f7f77777f7fafafffffafbfffff;

	lut_sub lut_578 ({sk[133], i_40_, i_22_, n_n834, n_n836, x415x, x423x}, x8563x);
	defparam lut_578.LUT_SIZE = 7;
	defparam lut_578.mask = 128'h77777f7f77777f7fffff8888fff08880;

	lut_sub lut_585 ({sk[134], i_40_, i_7_, i_32_, i_33_, x6939x}, n_n2581);
	defparam lut_585.LUT_SIZE = 6;
	defparam lut_585.mask = 64'h55ffffff10000000;

	lut_sub lut_587 ({sk[135], i_7_, i_39_, i_4_, i_36_, x81x, x80x}, n_n2838);
	defparam lut_587.LUT_SIZE = 7;
	defparam lut_587.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_589 ({sk[136], n_n1581, n_n1577, n_n1575, x7375x, x7382x}, x7386x);
	defparam lut_589.LUT_SIZE = 6;
	defparam lut_589.mask = 64'h55ffffff7fffffff;

	lut_sub lut_595 ({sk[137], n_n1908, x6958x, x6956x, x6957x, x8557x}, x7383x);
	defparam lut_595.LUT_SIZE = 6;
	defparam lut_595.mask = 64'h55ffffffbfffffff;

	lut_sub lut_601 ({sk[138], n_n560, x7432x, n_n1416, x696x, x1170x, x1171x}, n_n1409);
	defparam lut_601.LUT_SIZE = 7;
	defparam lut_601.mask = 128'h77777f7f77777f7f77ffffff7fffffff;

	lut_sub lut_607 ({sk[139], i_5_, i_12_, i_15_, x641x, x7391x, x7392x}, n_n1414);
	defparam lut_607.LUT_SIZE = 7;
	defparam lut_607.mask = 128'h77777f7f77777f7f7777777f77777777;

	lut_sub lut_611 ({sk[140], i_1_, i_2_, i_0_, x518x, x7402x, x8525x}, n_n1412);
	defparam lut_611.LUT_SIZE = 7;
	defparam lut_611.mask = 128'h77777f7f77777f7fbbbbbbbfbbbbbbbb;

	lut_sub lut_615 ({sk[141], i_39_, i_38_, i_37_, n_n459, x1187x, x7410x}, x7412x);
	defparam lut_615.LUT_SIZE = 7;
	defparam lut_615.mask = 128'h77777f7f77777f7f7f77777777777777;

	lut_sub lut_619 ({sk[142], x7440x, x7444x, x8523x, x8524x}, x7448x);
	defparam lut_619.LUT_SIZE = 5;
	defparam lut_619.mask = 32'h00ffefff;

	lut_sub lut_624 ({sk[143], i_23_, i_21_, n_n857, n_n860, n_n859, x40x}, x415x);
	defparam lut_624.LUT_SIZE = 7;
	defparam lut_624.mask = 128'h77777f7f77777f7f0007000000000000;

	lut_sub lut_627 ({sk[144], i_23_, i_21_, i_15_, i_19_, n_n857, x44x}, x423x);
	defparam lut_627.LUT_SIZE = 7;
	defparam lut_627.mask = 128'h77777f7f77777f7f0001000000000000;

	lut_sub lut_629 ({sk[145], n_n968, x82x, n_n960, x7455x, x132x, x475x}, n_n1651);
	defparam lut_629.LUT_SIZE = 7;
	defparam lut_629.mask = 128'h77777f7f77777f7f0f0f5f5f0f3f5f7f;

	lut_sub lut_633 ({sk[146], n_n969, n_n968, n_n1971, n_n1928, n_n819, x7462x}, x7463x);
	defparam lut_633.LUT_SIZE = 7;
	defparam lut_633.mask = 128'h77777f7f77777f7f5fff5fff5fff7fff;

	lut_sub lut_638 ({sk[147], i_15_, x313x, n_n833, x7478x, x1106x, x1104x}, n_n1484);
	defparam lut_638.LUT_SIZE = 7;
	defparam lut_638.mask = 128'h77777f7f77777f7f7f7f7fff5f5f5f5f;

	lut_sub lut_643 ({sk[148], x390x, x356x, x1073x, x1088x, x1089x, x7485x}, x7494x);
	defparam lut_643.LUT_SIZE = 7;
	defparam lut_643.mask = 128'h77777f7f77777f7f7fff7fff7fffffff;

	lut_sub lut_649 ({sk[149], i_12_, x362x, x428x, x691x, x1082x, x1074x}, x7495x);
	defparam lut_649.LUT_SIZE = 7;
	defparam lut_649.mask = 128'h77777f7f77777f7f7f7f7fff777777ff;

	lut_sub lut_654 ({sk[150], i_39_, i_15_, x392x, x791x, x1061x, x7497x}, n_n1489);
	defparam lut_654.LUT_SIZE = 7;
	defparam lut_654.mask = 128'h77777f7f77777f7f7fff77ff7f7f7777;

	lut_sub lut_659 ({sk[151], x335x, n_n685, x1049x, x1050x, x8521x, x8567x}, x7506x);
	defparam lut_659.LUT_SIZE = 7;
	defparam lut_659.mask = 128'h77777f7f77777f7fefffefffefffffff;

	lut_sub lut_665 ({sk[152], i_25_, n_n850, n_n848, x1044x, x1045x, x474x}, n_n1384);
	defparam lut_665.LUT_SIZE = 7;
	defparam lut_665.mask = 128'h77777f7f77777f7f0f0f0f0f0f3f0f7f;

	lut_sub lut_669 ({sk[153], i_39_, i_38_, i_37_}, n_n982);
	defparam lut_669.LUT_SIZE = 4;
	defparam lut_669.mask = 16'h1520;

	lut_sub lut_671 ({sk[154], i_7_, i_32_, i_34_, i_33_, i_36_, i_35_}, x328x);
	defparam lut_671.LUT_SIZE = 7;
	defparam lut_671.mask = 128'h77777f7f77777f7f0008000000000000;

	lut_sub lut_673 ({sk[155], i_40_, i_39_, i_38_, i_37_}, x325x);
	defparam lut_673.LUT_SIZE = 5;
	defparam lut_673.mask = 32'h00ff0008;

	lut_sub lut_675 ({sk[156], i_20_, i_21_, n_n411, x1038x, x486x, x303x}, x1031x);
	defparam lut_675.LUT_SIZE = 7;
	defparam lut_675.mask = 128'h77777f7f77777f7f0000000000000f1f;

	lut_sub lut_678 ({sk[157], i_25_, n_n853, n_n848, x532x, x474x}, x1032x);
	defparam lut_678.LUT_SIZE = 6;
	defparam lut_678.mask = 64'h55ffffff00003337;

	lut_sub lut_681 ({sk[158], o_15_, x84x, x347x, x407x, x7524x, x8520x}, x7530x);
	defparam lut_681.LUT_SIZE = 7;
	defparam lut_681.mask = 128'h77777f7f77777f7fbbbbbbbfffffffff;

	lut_sub lut_686 ({sk[159], i_12_, i_11_, i_17_, i_16_, i_15_, x317x}, x109x);
	defparam lut_686.LUT_SIZE = 7;
	defparam lut_686.mask = 128'h77777f7f77777f7f0000010101110000;

	lut_sub lut_690 ({sk[160], i_12_, i_11_, x478x, n_n1048, n_n785, x407x}, n_n1372);
	defparam lut_690.LUT_SIZE = 7;
	defparam lut_690.mask = 128'h77777f7f77777f7f0003010301030003;

	lut_sub lut_694 ({sk[161], i_32_, i_31_, i_33_}, n_n1048);
	defparam lut_694.LUT_SIZE = 4;
	defparam lut_694.mask = 16'h1540;

	lut_sub lut_696 ({sk[162], i_40_, i_34_, i_36_, i_35_, i_37_, n_n960}, n_n785);
	defparam lut_696.LUT_SIZE = 7;
	defparam lut_696.mask = 128'h77777f7f77777f7f0000000040000000;

	lut_sub lut_698 ({sk[163], i_17_, i_16_, n_n775, n_n1048, x98x, x522x}, x7526x);
	defparam lut_698.LUT_SIZE = 7;
	defparam lut_698.mask = 128'h77777f7f77777f7f0000000700070007;

	lut_sub lut_703 ({sk[164], i_23_, i_15_, x359x, x57x, n_n1023, n_n428}, n_n1375);
	defparam lut_703.LUT_SIZE = 7;
	defparam lut_703.mask = 128'h77777f7f77777f7f0000000000000001;

	lut_sub lut_705 ({sk[165], i_19_, x359x, n_n1023, x484x, x380x, x7124x}, n_n1374);
	defparam lut_705.LUT_SIZE = 7;
	defparam lut_705.mask = 128'h77777f7f77777f7f0000000000000015;

	lut_sub lut_708 ({sk[166], x122x, x7535x, x7536x, x7537x, x8519x}, n_n1356);
	defparam lut_708.LUT_SIZE = 6;
	defparam lut_708.mask = 64'h55ffffffbfffffff;

	lut_sub lut_714 ({sk[167], n_n1373, n_n949, x480x, x386x, x997x, x998x}, x7546x);
	defparam lut_714.LUT_SIZE = 7;
	defparam lut_714.mask = 128'h77777f7f77777f7f7777777fffffffff;

	lut_sub lut_719 ({sk[168], i_22_, x247x, x99x, n_n1072, x417x, x380x}, x7547x);
	defparam lut_719.LUT_SIZE = 7;
	defparam lut_719.mask = 128'h77777f7f77777f7f0303ffff0307ffff;

	lut_sub lut_723 ({sk[169], i_40_, i_39_}, n_n1064);
	defparam lut_723.LUT_SIZE = 3;
	defparam lut_723.mask = 8'h32;

	lut_sub lut_725 ({sk[170], i_40_, i_39_, i_12_, i_11_, x45x, n_n693}, x146x);
	defparam lut_725.LUT_SIZE = 7;
	defparam lut_725.mask = 128'h77777f7f77777f7f0000000000000010;

	lut_sub lut_727 ({sk[171], i_32_, i_34_, i_33_, i_36_, i_35_, i_37_}, x340x);
	defparam lut_727.LUT_SIZE = 7;
	defparam lut_727.mask = 128'h77777f7f77777f7f0000004000000000;

	lut_sub lut_729 ({sk[172], x7621x, x7622x, x7636x, x7637x, x8554x}, x7639x);
	defparam lut_729.LUT_SIZE = 6;
	defparam lut_729.mask = 64'h55ffffffbfffffff;

	lut_sub lut_735 ({sk[173], n_n1283, n_n1285, x7591x, x7614x}, x7616x);
	defparam lut_735.LUT_SIZE = 5;
	defparam lut_735.mask = 32'h00ff7fff;

	lut_sub lut_740 ({sk[174], n_n833, n_n837, n_n834, x7560x, x8559x}, n_n1280);
	defparam lut_740.LUT_SIZE = 6;
	defparam lut_740.mask = 64'h55ffffffbbbbbfff;

	lut_sub lut_745 ({sk[175], i_40_, x148x, x7565x, x7566x, x7567x, x7568x}, n_n1282);
	defparam lut_745.LUT_SIZE = 7;
	defparam lut_745.mask = 128'h77777f7f77777f7f7fff7fff7fffffff;

	lut_sub lut_751 ({sk[176], x329x, n_n926, n_n764, x365x, x395x, x962x}, x7574x);
	defparam lut_751.LUT_SIZE = 7;
	defparam lut_751.mask = 128'h77777f7f77777f7f575757ff777777ff;

	lut_sub lut_756 ({sk[177], x7605x, x912x, x913x, x927x, x7604x}, x7615x);
	defparam lut_756.LUT_SIZE = 6;
	defparam lut_756.mask = 64'h55ffffff7fffffff;

	lut_sub lut_762 ({sk[178], n_n1330, n_n1332, n_n1326, x7660x, x7681x}, x7684x);
	defparam lut_762.LUT_SIZE = 6;
	defparam lut_762.mask = 64'h55ffffff7fffffff;

	lut_sub lut_768 ({sk[179], i_40_, n_n795, x358x, x100x, n_n710, x756x}, x536x);
	defparam lut_768.LUT_SIZE = 7;
	defparam lut_768.mask = 128'h77777f7f77777f7f0003555700000000;

	lut_sub lut_771 ({sk[180], i_40_, n_n985, n_n525, x854x, x7667x, x8516x}, n_n1329);
	defparam lut_771.LUT_SIZE = 7;
	defparam lut_771.mask = 128'h77777f7f77777f7fbbbbbfbfbbbbbfff;

	lut_sub lut_776 ({sk[181], x7663x, x519x, x858x, x7662x, x7672x}, x7674x);
	defparam lut_776.LUT_SIZE = 6;
	defparam lut_776.mask = 64'h55ffffff7fffffff;

	lut_sub lut_782 ({sk[182], i_15_, x287x, x282x, x283x, x289x, x7720x}, x7732x);
	defparam lut_782.LUT_SIZE = 7;
	defparam lut_782.mask = 128'h77777f7f77777f7f7777ffff7fffffff;

	lut_sub lut_788 ({sk[183], n_n1203, x7733x, x7735x, x7737x, x8514x}, n_n1184);
	defparam lut_788.LUT_SIZE = 6;
	defparam lut_788.mask = 64'h55ffffffbfffffff;

	lut_sub lut_794 ({sk[184], x45x, x517x, x7713x, n_n918, x7714x, x7715x}, n_n1197);
	defparam lut_794.LUT_SIZE = 7;
	defparam lut_794.mask = 128'h77777f7f77777f7f7777777777ff7fff;

	lut_sub lut_799 ({sk[185], i_32_, n_n926, n_n1066, x513x, x275x, x7729x}, x7730x);
	defparam lut_799.LUT_SIZE = 7;
	defparam lut_799.mask = 128'h77777f7f77777f7f7777777f77777777;

	lut_sub lut_803 ({sk[186], i_2_, x384x, x249x, x216x, x7746x, x8513x}, x7763x);
	defparam lut_803.LUT_SIZE = 7;
	defparam lut_803.mask = 128'h77777f7f77777f7fbfffbfffbfffffff;

	lut_sub lut_809 ({sk[187], n_n1195, n_n1193, x311x, x7702x, x7703x, x7762x}, x7764x);
	defparam lut_809.LUT_SIZE = 7;
	defparam lut_809.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_816 ({sk[188], x7793x, n_n1235, x7814x, n_n1242, n_n1237, n_n1239}, x7824x);
	defparam lut_816.LUT_SIZE = 7;
	defparam lut_816.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_823 ({sk[189], i_14_, i_12_, i_15_, n_n860, n_n642, x114x}, x483x);
	defparam lut_823.LUT_SIZE = 7;
	defparam lut_823.mask = 128'h77777f7f77777f7f0011001300110011;

	lut_sub lut_826 ({sk[190], i_12_, i_11_, i_15_, n_n860, x38x, x126x}, x7820x);
	defparam lut_826.LUT_SIZE = 7;
	defparam lut_826.mask = 128'h77777f7f77777f7f0505050705070505;

	lut_sub lut_830 ({sk[191], i_14_, i_17_, i_16_, i_32_, i_33_, x87x}, x463x);
	defparam lut_830.LUT_SIZE = 7;
	defparam lut_830.mask = 128'h77777f7f77777f7f0000001000000000;

	lut_sub lut_832 ({sk[192], i_12_, n_n775, x341x, n_n860, x483x, x7820x}, x7821x);
	defparam lut_832.LUT_SIZE = 7;
	defparam lut_832.mask = 128'h77777f7f77777f7f00007777000f777f;

	lut_sub lut_836 ({sk[193], i_14_, n_n1074, n_n560, x407x, x39x, x686x}, x1923x);
	defparam lut_836.LUT_SIZE = 7;
	defparam lut_836.mask = 128'h77777f7f77777f7f0000005700000003;

	lut_sub lut_839 ({sk[194], i_17_, i_16_, x45x, x92x, x36x, x484x}, x6726x);
	defparam lut_839.LUT_SIZE = 7;
	defparam lut_839.mask = 128'h77777f7f77777f7f0000000500050007;

	lut_sub lut_843 ({sk[195], i_40_, i_7_, i_39_, i_33_, i_38_, x503x}, x145x);
	defparam lut_843.LUT_SIZE = 7;
	defparam lut_843.mask = 128'h77777f7f77777f7f00000f0f11001f0f;

	lut_sub lut_846 ({sk[196], i_17_, i_16_, n_n1074, n_n560, x98x, x522x}, x1883x);
	defparam lut_846.LUT_SIZE = 7;
	defparam lut_846.mask = 128'h77777f7f77777f7f0000000700070007;

	lut_sub lut_851 ({sk[197], i_26_, n_n709, n_n1015, x324x, x391x, n_n1021}, x6752x);
	defparam lut_851.LUT_SIZE = 7;
	defparam lut_851.mask = 128'h77777f7f77777f7f1133113311331f3f;

	lut_sub lut_855 ({sk[198], i_36_, i_38_, i_37_}, n_n985);
	defparam lut_855.LUT_SIZE = 4;
	defparam lut_855.mask = 16'h1540;

	lut_sub lut_857 ({sk[199], i_7_, i_3_, i_4_, i_1_, i_2_, x80x}, n_n515);
	defparam lut_857.LUT_SIZE = 7;
	defparam lut_857.mask = 128'h77777f7f77777f7f4000000000000000;

	lut_sub lut_859 ({sk[200], i_40_, i_39_}, n_n1008);
	defparam lut_859.LUT_SIZE = 3;
	defparam lut_859.mask = 8'h38;

	lut_sub lut_861 ({sk[201], n_n1011, n_n842, n_n1067, x335x, x373x, x89x}, x1867x);
	defparam lut_861.LUT_SIZE = 7;
	defparam lut_861.mask = 128'h77777f7f77777f7f0000001f0000005f;

	lut_sub lut_865 ({sk[202], i_40_, n_n979, n_n982, n_n861, n_n795, x358x}, x6767x);
	defparam lut_865.LUT_SIZE = 7;
	defparam lut_865.mask = 128'h77777f7f77777f7f0000000f11111111;

	lut_sub lut_868 ({sk[203], i_39_, i_38_, i_37_, x88x, n_n991, x528x}, x6768x);
	defparam lut_868.LUT_SIZE = 7;
	defparam lut_868.mask = 128'h77777f7f77777f7f0003000055000000;

	lut_sub lut_871 ({sk[204], i_4_, i_1_, x314x, x6818x, n_n926, x6813x}, n_n1083);
	defparam lut_871.LUT_SIZE = 7;
	defparam lut_871.mask = 128'h77777f7f77777f7f5f5f5f7f5f7f5f7f;

	lut_sub lut_876 ({sk[205], n_n709, n_n287, x238x, x1805x, x6829x, x6830x}, n_n1084);
	defparam lut_876.LUT_SIZE = 7;
	defparam lut_876.mask = 128'h77777f7f77777f7f7fff7fff7fffffff;

	lut_sub lut_882 ({sk[206], i_7_, i_1_, i_2_, i_0_, n_n1074, x95x}, x1706x);
	defparam lut_882.LUT_SIZE = 7;
	defparam lut_882.mask = 128'h77777f7f77777f7f0101000100000000;

	lut_sub lut_885 ({sk[207], i_40_, i_39_, i_38_, n_n330, x51x, x328x}, x6922x);
	defparam lut_885.LUT_SIZE = 7;
	defparam lut_885.mask = 128'h77777f7f77777f7f0300000000550000;

	lut_sub lut_888 ({sk[208], n_n978, n_n998, n_n973, n_n158, x35x, x385x}, x6923x);
	defparam lut_888.LUT_SIZE = 7;
	defparam lut_888.mask = 128'h77777f7f77777f7f0000000355555557;

	lut_sub lut_891 ({sk[209], n_n1021, x93x, x6819x, x6820x, x313x, x6920x}, x8544x);
	defparam lut_891.LUT_SIZE = 7;
	defparam lut_891.mask = 128'h77777f7f77777f7ffffff000eeeee000;

	lut_sub lut_898 ({sk[210], i_7_, i_5_, i_12_, i_11_}, x35x);
	defparam lut_898.LUT_SIZE = 5;
	defparam lut_898.mask = 32'h00ff7000;

	lut_sub lut_901 ({sk[211], i_40_, i_39_, i_38_, n_n964, x76x, x6862x}, n_n1936);
	defparam lut_901.LUT_SIZE = 7;
	defparam lut_901.mask = 128'h77777f7f77777f7f0000000000010000;

	lut_sub lut_903 ({sk[212], i_22_, i_38_, n_n1014, x52x, x340x, x304x}, x552x);
	defparam lut_903.LUT_SIZE = 7;
	defparam lut_903.mask = 128'h77777f7f77777f7f0505050505370505;

	lut_sub lut_906 ({sk[213], i_21_, i_15_, n_n853, n_n850, n_n469, x52x}, x1694x);
	defparam lut_906.LUT_SIZE = 7;
	defparam lut_906.mask = 128'h77777f7f77777f7f0000011100000000;

	lut_sub lut_909 ({sk[214], i_32_, i_33_}, x46x);
	defparam lut_909.LUT_SIZE = 3;
	defparam lut_909.mask = 8'h34;

	lut_sub lut_911 ({sk[215], i_7_, i_2_, i_0_, i_32_, i_34_, i_33_}, x429x);
	defparam lut_911.LUT_SIZE = 7;
	defparam lut_911.mask = 128'h77777f7f77777f7f0000004000000000;

	lut_sub lut_913 ({sk[216], i_7_, i_39_, i_1_, i_36_, x81x, x80x}, n_n2836);
	defparam lut_913.LUT_SIZE = 7;
	defparam lut_913.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_915 ({sk[217], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x71x);
	defparam lut_915.LUT_SIZE = 7;
	defparam lut_915.mask = 128'h77777f7f77777f7f0004000000100020;

	lut_sub lut_919 ({sk[218], i_7_, i_3_, i_0_, i_32_, i_34_, i_33_}, x302x);
	defparam lut_919.LUT_SIZE = 7;
	defparam lut_919.mask = 128'h77777f7f77777f7f0000004000000000;

	lut_sub lut_921 ({sk[219], i_4_, n_n2581, x431x, x541x, x350x, x362x}, x8540x);
	defparam lut_921.LUT_SIZE = 7;
	defparam lut_921.mask = 128'h77777f7f77777f7ffaf00000eae00000;

	lut_sub lut_926 ({sk[220], i_39_, i_36_, i_38_, i_37_}, n_n926);
	defparam lut_926.LUT_SIZE = 5;
	defparam lut_926.mask = 32'h00ff4000;

	lut_sub lut_928 ({sk[221], i_40_, i_39_, i_36_, i_38_, i_37_}, x92x);
	defparam lut_928.LUT_SIZE = 6;
	defparam lut_928.mask = 64'h55ffffff00000020;

	lut_sub lut_930 ({sk[222], i_16_, i_34_, i_33_, i_35_, n_n933}, x319x);
	defparam lut_930.LUT_SIZE = 6;
	defparam lut_930.mask = 64'h55ffffff00000400;

	lut_sub lut_932 ({sk[223], i_7_, i_5_, i_12_, i_11_, i_15_}, x470x);
	defparam lut_932.LUT_SIZE = 6;
	defparam lut_932.mask = 64'h55ffffff10000000;

	lut_sub lut_934 ({sk[224], i_16_, x425x, x78x, n_n527, x388x, x7015x}, x7018x);
	defparam lut_934.LUT_SIZE = 7;
	defparam lut_934.mask = 128'h77777f7f77777f7f111155551111555f;

	lut_sub lut_938 ({sk[225], i_31_, i_35_, x46x, n_n462, x7019x, x7020x}, x7021x);
	defparam lut_938.LUT_SIZE = 7;
	defparam lut_938.mask = 128'h77777f7f77777f7f5557555555555555;

	lut_sub lut_941 ({sk[226], i_40_, i_7_, i_32_, i_33_}, x88x);
	defparam lut_941.LUT_SIZE = 5;
	defparam lut_941.mask = 32'h00ff4000;

	lut_sub lut_943 ({sk[227], n_n1074, n_n880, x326x, x490x, n_n700, x7235x}, x7237x);
	defparam lut_943.LUT_SIZE = 7;
	defparam lut_943.mask = 128'h77777f7f77777f7f55555757555557ff;

	lut_sub lut_947 ({sk[228], i_2_, i_38_, i_37_, x77x, x464x, x7259x}, x7261x);
	defparam lut_947.LUT_SIZE = 7;
	defparam lut_947.mask = 128'h77777f7f77777f7f57575555575f5555;

	lut_sub lut_951 ({sk[229], i_0_, i_38_, n_n700, n_n1073, x397x, x1361x}, x1356x);
	defparam lut_951.LUT_SIZE = 7;
	defparam lut_951.mask = 128'h77777f7f77777f7f0000555f0000777f;

	lut_sub lut_955 ({sk[230], i_9_, i_39_, i_16_, i_36_, x45x, x1333x}, x7260x);
	defparam lut_955.LUT_SIZE = 7;
	defparam lut_955.mask = 128'h77777f7f77777f7f5555755555555555;

	lut_sub lut_958 ({sk[231], i_39_, i_38_, x90x, x46x, x389x, x810x}, x8531x);
	defparam lut_958.LUT_SIZE = 7;
	defparam lut_958.mask = 128'h77777f7f77777f7ffa00fafac800c8c8;

	lut_sub lut_967 ({sk[232], i_40_, n_n688, n_n918, x726x, x725x, x1266x}, x7329x);
	defparam lut_967.LUT_SIZE = 7;
	defparam lut_967.mask = 128'h77777f7f77777f7f55555f5f55775577;

	lut_sub lut_971 ({sk[233], x313x, x6920x, x85x, x7339x, x1245x, x7340x}, n_n1447);
	defparam lut_971.LUT_SIZE = 7;
	defparam lut_971.mask = 128'h77777f7f77777f7f777f777f777fffff;

	lut_sub lut_976 ({sk[234], n_n559, x130x, x327x, n_n550, x139x, x1277x}, n_n1453);
	defparam lut_976.LUT_SIZE = 7;
	defparam lut_976.mask = 128'h77777f7f77777f7f555fffff777fffff;

	lut_sub lut_981 ({sk[235], n_n560, x364x, x336x, n_n550, x7321x, x7319x}, n_n1452);
	defparam lut_981.LUT_SIZE = 7;
	defparam lut_981.mask = 128'h77777f7f77777f7f777777ff7f7f7fff;

	lut_sub lut_986 ({sk[236], x528x, x100x, x1254x, x7335x, x7336x, x7343x}, x7344x);
	defparam lut_986.LUT_SIZE = 7;
	defparam lut_986.mask = 128'h77777f7f77777f7f7fff7fff7fffffff;

	lut_sub lut_992 ({sk[237], i_39_, i_36_, i_35_, i_38_, i_37_}, n_n560);
	defparam lut_992.LUT_SIZE = 6;
	defparam lut_992.mask = 64'h55ffffff40000000;

	lut_sub lut_994 ({sk[238], x338x, x60x, x7406x, x1161x, x1163x, x7429x}, x7432x);
	defparam lut_994.LUT_SIZE = 7;
	defparam lut_994.mask = 128'h77777f7f77777f7f7f7f7f7f7f7f7fff;

	lut_sub lut_999 ({sk[239], x76x, x517x, x103x, x1179x, x1181x, x7417x}, n_n1416);
	defparam lut_999.LUT_SIZE = 7;
	defparam lut_999.mask = 128'h77777f7f77777f7f7f7f7f7f7f7f7fff;

	lut_sub lut_1004 ({sk[240], i_17_, i_16_, i_15_, n_n488, x76x, x7426x}, x696x);
	defparam lut_1004.LUT_SIZE = 7;
	defparam lut_1004.mask = 128'h77777f7f77777f7f5557555755575555;

	lut_sub lut_1008 ({sk[241], i_17_, i_16_, i_31_, n_n1074, x36x, x327x}, x1170x);
	defparam lut_1008.LUT_SIZE = 7;
	defparam lut_1008.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_1010 ({sk[242], n_n1073, n_n492, n_n488, x76x, x352x, x343x}, x1171x);
	defparam lut_1010.LUT_SIZE = 7;
	defparam lut_1010.mask = 128'h77777f7f77777f7f0000000000010101;

	lut_sub lut_1013 ({sk[243], i_39_, i_36_, i_38_, i_37_}, n_n833);
	defparam lut_1013.LUT_SIZE = 5;
	defparam lut_1013.mask = 32'h00ff0020;

	lut_sub lut_1015 ({sk[244], i_7_, i_32_, i_31_, n_n1066, x718x, x7477x}, x7478x);
	defparam lut_1015.LUT_SIZE = 7;
	defparam lut_1015.mask = 128'h77777f7f77777f7f5557555555555555;

	lut_sub lut_1018 ({sk[245], i_40_, n_n795, n_n976, x376x, x1109x, x1110x}, x1106x);
	defparam lut_1018.LUT_SIZE = 7;
	defparam lut_1018.mask = 128'h77777f7f77777f7f000000003737373f;

	lut_sub lut_1022 ({sk[246], i_39_, i_36_, i_38_, i_37_, n_n1066, n_n668}, x1104x);
	defparam lut_1022.LUT_SIZE = 7;
	defparam lut_1022.mask = 128'h77777f7f77777f7f1011000011010000;

	lut_sub lut_1027 ({sk[247], i_7_, i_5_, i_12_}, n_n850);
	defparam lut_1027.LUT_SIZE = 4;
	defparam lut_1027.mask = 16'h1540;

	lut_sub lut_1029 ({sk[248], i_21_, i_22_, i_15_}, n_n848);
	defparam lut_1029.LUT_SIZE = 4;
	defparam lut_1029.mask = 16'h1501;

	lut_sub lut_1031 ({sk[249], i_40_, i_20_, i_39_, i_38_, x364x, x77x}, x1044x);
	defparam lut_1031.LUT_SIZE = 7;
	defparam lut_1031.mask = 128'h77777f7f77777f7f0000000000000010;

	lut_sub lut_1033 ({sk[250], i_24_, n_n853, n_n850, x50x, x101x, x1047x}, x1045x);
	defparam lut_1033.LUT_SIZE = 7;
	defparam lut_1033.mask = 128'h77777f7f77777f7f0000000000575757;

	lut_sub lut_1038 ({sk[251], i_39_, i_23_, i_24_, i_38_, n_n1074, n_n968}, x474x);
	defparam lut_1038.LUT_SIZE = 7;
	defparam lut_1038.mask = 128'h77777f7f77777f7f0000000000000001;

	lut_sub lut_1040 ({sk[252], i_32_, i_31_, i_33_, i_37_, n_n1011, n_n1047}, x84x);
	defparam lut_1040.LUT_SIZE = 7;
	defparam lut_1040.mask = 128'h77777f7f77777f7f0001000000000000;

	lut_sub lut_1042 ({sk[253], i_12_, i_11_}, x347x);
	defparam lut_1042.LUT_SIZE = 3;
	defparam lut_1042.mask = 8'h32;

	lut_sub lut_1044 ({sk[254], i_5_, i_17_, i_16_, i_15_}, x407x);
	defparam lut_1044.LUT_SIZE = 5;
	defparam lut_1044.mask = 32'h00ff0100;

	lut_sub lut_1046 ({sk[255], i_28_, i_29_, n_n2687, x361x, x457x}, x7524x);
	defparam lut_1046.LUT_SIZE = 6;
	defparam lut_1046.mask = 64'h55ffffff1f0f0f0f;

	lut_sub lut_1049 ({sk[256], i_19_, x48x, x72x, n_n411, n_n857, x57x}, x8520x);
	defparam lut_1049.LUT_SIZE = 7;
	defparam lut_1049.mask = 128'h77777f7f77777f7ffffffefefffcfefc;

	lut_sub lut_1056 ({sk[257], i_40_, i_7_, i_12_, i_32_, x525x, x8568x}, x7621x);
	defparam lut_1056.LUT_SIZE = 7;
	defparam lut_1056.mask = 128'h77777f7f77777f7f00300000aabaaaaa;

	lut_sub lut_1059 ({sk[258], i_40_, i_7_, x46x, n_n982, n_n998, n_n2836}, x7622x);
	defparam lut_1059.LUT_SIZE = 7;
	defparam lut_1059.mask = 128'h77777f7f77777f7f5557555555555555;

	lut_sub lut_1062 ({sk[259], x7555x, x986x, x7552x, x7553x, x7634x}, x7636x);
	defparam lut_1062.LUT_SIZE = 6;
	defparam lut_1062.mask = 64'h55ffffff7fffffff;

	lut_sub lut_1068 ({sk[260], i_37_, n_n1014, x328x, x131x, x891x, x892x}, x7637x);
	defparam lut_1068.LUT_SIZE = 7;
	defparam lut_1068.mask = 128'h77777f7f77777f7f7f7f7fff7f7f7f7f;

	lut_sub lut_1073 ({sk[261], i_7_, i_3_, i_4_, i_1_, n_n833, x80x}, x8554x);
	defparam lut_1073.LUT_SIZE = 7;
	defparam lut_1073.mask = 128'h77777f7f77777f7ffeeeeeeeffffffff;

	lut_sub lut_1078 ({sk[262], i_31_, x45x, x506x, x882x, x883x, x884x}, n_n1330);
	defparam lut_1078.LUT_SIZE = 7;
	defparam lut_1078.mask = 128'h77777f7f77777f7f7f7f7fff7f7f7f7f;

	lut_sub lut_1083 ({sk[263], x878x, x130x, x877x}, n_n1332);
	defparam lut_1083.LUT_SIZE = 4;
	defparam lut_1083.mask = 16'h157f;

	lut_sub lut_1087 ({sk[264], x358x, n_n977, n_n710, x7655x, x870x, x7653x}, n_n1326);
	defparam lut_1087.LUT_SIZE = 7;
	defparam lut_1087.mask = 128'h77777f7f77777f7f7f7f7f7f7f7f7fff;

	lut_sub lut_1092 ({sk[265], n_n795, x435x, x131x, x499x, x177x, x7657x}, x7660x);
	defparam lut_1092.LUT_SIZE = 7;
	defparam lut_1092.mask = 128'h77777f7f77777f7f77ff77ff7fffffff;

	lut_sub lut_1098 ({sk[266], x316x, x94x, x507x, x106x, x466x, x477x}, x7681x);
	defparam lut_1098.LUT_SIZE = 7;
	defparam lut_1098.mask = 128'h77777f7f77777f7f7777777777ff7fff;

	lut_sub lut_1103 ({sk[267], x358x, n_n883, n_n710, x189x, x7789x, x7790x}, x7793x);
	defparam lut_1103.LUT_SIZE = 7;
	defparam lut_1103.mask = 128'h77777f7f77777f7f7f7f7f7f7f7f7fff;

	lut_sub lut_1108 ({sk[268], i_39_, i_26_, x439x, x168x, x7798x, x7799x}, n_n1235);
	defparam lut_1108.LUT_SIZE = 7;
	defparam lut_1108.mask = 128'h77777f7f77777f7f7fff7f7f7f7f7f7f;

	lut_sub lut_1113 ({sk[269], i_15_, x47x, x339x, x147x, x7810x, x7812x}, x7814x);
	defparam lut_1113.LUT_SIZE = 7;
	defparam lut_1113.mask = 128'h77777f7f77777f7f7f7f7fff7f7f7f7f;

	lut_sub lut_1118 ({sk[270], i_23_, i_37_, n_n880, x129x, x136x, x137x}, n_n1242);
	defparam lut_1118.LUT_SIZE = 7;
	defparam lut_1118.mask = 128'h77777f7f77777f7f0f0f0f0f0f0f0f7f;

	lut_sub lut_1122 ({sk[271], i_39_, i_25_, x7775x, x439x, x212x, x7773x}, n_n1237);
	defparam lut_1122.LUT_SIZE = 7;
	defparam lut_1122.mask = 128'h77777f7f77777f7f77ff7fff77ff77ff;

	lut_sub lut_1127 ({sk[272], i_40_, x663x, x7784x, x7785x, x7786x}, n_n1239);
	defparam lut_1127.LUT_SIZE = 6;
	defparam lut_1127.mask = 64'h55ffffff7f7f7fff;

	lut_sub lut_1132 ({sk[273], i_9_, i_5_}, x317x);
	defparam lut_1132.LUT_SIZE = 3;
	defparam lut_1132.mask = 8'h32;

	lut_sub lut_1134 ({sk[274], i_9_, i_5_, i_11_}, n_n955);
	defparam lut_1134.LUT_SIZE = 4;
	defparam lut_1134.mask = 16'h1504;

	lut_sub lut_1136 ({sk[275], i_34_, i_36_, i_35_}, n_n1047);
	defparam lut_1136.LUT_SIZE = 4;
	defparam lut_1136.mask = 16'h1580;

	lut_sub lut_1138 ({sk[276], i_5_, i_13_, i_12_, i_11_, i_32_, i_33_}, x399x);
	defparam lut_1138.LUT_SIZE = 7;
	defparam lut_1138.mask = 128'h77777f7f77777f7f4000000000000000;

	lut_sub lut_1140 ({sk[277], i_40_, i_39_, i_38_, i_37_, n_n1047, x399x}, x1934x);
	defparam lut_1140.LUT_SIZE = 7;
	defparam lut_1140.mask = 128'h77777f7f77777f7f0100100011001010;

	lut_sub lut_1145 ({sk[278], i_38_, i_37_}, n_n709);
	defparam lut_1145.LUT_SIZE = 3;
	defparam lut_1145.mask = 8'h38;

	lut_sub lut_1147 ({sk[279], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x327x);
	defparam lut_1147.LUT_SIZE = 7;
	defparam lut_1147.mask = 128'h77777f7f77777f7f0000000000002000;

	lut_sub lut_1149 ({sk[280], i_9_, i_17_, i_16_, i_15_, x327x}, x6722x);
	defparam lut_1149.LUT_SIZE = 6;
	defparam lut_1149.mask = 64'h55ffffff00010111;

	lut_sub lut_1153 ({sk[281], i_32_, i_34_, i_33_}, n_n1074);
	defparam lut_1153.LUT_SIZE = 4;
	defparam lut_1153.mask = 16'h1540;

	lut_sub lut_1155 ({sk[282], i_14_, i_12_, i_11_, x6722x, n_n1074}, n_n1159);
	defparam lut_1155.LUT_SIZE = 6;
	defparam lut_1155.mask = 64'h55ffffff00000001;

	lut_sub lut_1157 ({sk[283], i_12_, i_11_}, x39x);
	defparam lut_1157.LUT_SIZE = 3;
	defparam lut_1157.mask = 8'h36;

	lut_sub lut_1160 ({sk[284], i_9_, i_5_, i_12_, i_17_, i_16_, i_15_}, x686x);
	defparam lut_1160.LUT_SIZE = 7;
	defparam lut_1160.mask = 128'h77777f7f77777f7f0001000000150000;

	lut_sub lut_1164 ({sk[285], i_32_, i_34_, i_33_, i_35_}, x45x);
	defparam lut_1164.LUT_SIZE = 5;
	defparam lut_1164.mask = 32'h00ff2000;

	lut_sub lut_1166 ({sk[286], i_5_, i_12_, i_11_, i_15_}, x36x);
	defparam lut_1166.LUT_SIZE = 5;
	defparam lut_1166.mask = 32'h00ff1500;

	lut_sub lut_1169 ({sk[287], i_9_, i_5_, i_12_, i_15_}, x484x);
	defparam lut_1169.LUT_SIZE = 5;
	defparam lut_1169.mask = 32'h00ff0010;

	lut_sub lut_1171 ({sk[288], i_40_, i_34_, i_33_, i_36_, n_n990}, x525x);
	defparam lut_1171.LUT_SIZE = 6;
	defparam lut_1171.mask = 64'h55ffffff00000100;

	lut_sub lut_1173 ({sk[289], x90x, n_n880, n_n874, x357x, n_n884, x233x}, x1913x);
	defparam lut_1173.LUT_SIZE = 7;
	defparam lut_1173.mask = 128'h77777f7f77777f7f1113111311133333;

	lut_sub lut_1177 ({sk[290], i_5_, i_31_, x46x, n_n1047, x55x, x331x}, x1912x);
	defparam lut_1177.LUT_SIZE = 7;
	defparam lut_1177.mask = 128'h77777f7f77777f7f0000555700000000;

	lut_sub lut_1180 ({sk[291], i_9_, i_5_, i_16_, x389x, x339x, n_n1072}, x6733x);
	defparam lut_1180.LUT_SIZE = 7;
	defparam lut_1180.mask = 128'h77777f7f77777f7f3705050505050505;

	lut_sub lut_1183 ({sk[292], i_39_, i_38_}, n_n1015);
	defparam lut_1183.LUT_SIZE = 3;
	defparam lut_1183.mask = 8'h32;

	lut_sub lut_1185 ({sk[293], i_40_, i_39_, i_38_}, x66x);
	defparam lut_1185.LUT_SIZE = 4;
	defparam lut_1185.mask = 16'h1523;

	lut_sub lut_1188 ({sk[294], i_32_, i_34_, i_33_, i_36_, i_35_, i_37_}, x90x);
	defparam lut_1188.LUT_SIZE = 7;
	defparam lut_1188.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_1190 ({sk[295], i_32_, i_34_, i_33_, i_35_, i_37_}, x503x);
	defparam lut_1190.LUT_SIZE = 6;
	defparam lut_1190.mask = 64'h55ffffff02000000;

	lut_sub lut_1192 ({sk[296], i_34_, i_36_, i_35_}, n_n1002);
	defparam lut_1192.LUT_SIZE = 4;
	defparam lut_1192.mask = 16'h1510;

	lut_sub lut_1194 ({sk[297], i_32_, i_34_, i_33_, i_36_, i_35_}, x324x);
	defparam lut_1194.LUT_SIZE = 6;
	defparam lut_1194.mask = 64'h55ffffff01000000;

	lut_sub lut_1196 ({sk[298], i_36_, i_35_, i_37_}, n_n864);
	defparam lut_1196.LUT_SIZE = 4;
	defparam lut_1196.mask = 16'h1502;

	lut_sub lut_1198 ({sk[299], i_34_, i_33_, i_35_}, n_n1066);
	defparam lut_1198.LUT_SIZE = 4;
	defparam lut_1198.mask = 16'h1520;

	lut_sub lut_1200 ({sk[300], i_17_, i_16_, i_32_, n_n1014, n_n1009, n_n1066}, x537x);
	defparam lut_1200.LUT_SIZE = 7;
	defparam lut_1200.mask = 128'h77777f7f77777f7f0000010001000100;

	lut_sub lut_1203 ({sk[301], i_9_, i_5_, i_12_, i_11_, i_17_, i_15_}, x478x);
	defparam lut_1203.LUT_SIZE = 7;
	defparam lut_1203.mask = 128'h77777f7f77777f7f0000000001000000;

	lut_sub lut_1205 ({sk[302], i_40_, i_39_}, n_n1021);
	defparam lut_1205.LUT_SIZE = 3;
	defparam lut_1205.mask = 8'h34;

	lut_sub lut_1207 ({sk[303], i_39_, i_38_, i_37_}, n_n1055);
	defparam lut_1207.LUT_SIZE = 4;
	defparam lut_1207.mask = 16'h1540;

	lut_sub lut_1209 ({sk[304], i_38_, i_37_}, x81x);
	defparam lut_1209.LUT_SIZE = 3;
	defparam lut_1209.mask = 8'h34;

	lut_sub lut_1211 ({sk[305], i_7_, i_32_, i_34_, i_33_, i_35_}, x314x);
	defparam lut_1211.LUT_SIZE = 6;
	defparam lut_1211.mask = 64'h55ffffff02000000;

	lut_sub lut_1213 ({sk[306], i_32_, i_34_, i_33_, i_35_}, x80x);
	defparam lut_1213.LUT_SIZE = 5;
	defparam lut_1213.mask = 32'h00ff0200;

	lut_sub lut_1215 ({sk[307], i_7_, i_3_, i_4_}, n_n842);
	defparam lut_1215.LUT_SIZE = 4;
	defparam lut_1215.mask = 16'h1540;

	lut_sub lut_1217 ({sk[308], i_1_, i_2_, i_0_}, n_n1067);
	defparam lut_1217.LUT_SIZE = 4;
	defparam lut_1217.mask = 16'h1540;

	lut_sub lut_1219 ({sk[309], i_38_, i_37_}, x316x);
	defparam lut_1219.LUT_SIZE = 3;
	defparam lut_1219.mask = 8'h32;

	lut_sub lut_1221 ({sk[310], i_39_, i_38_, i_37_}, n_n990);
	defparam lut_1221.LUT_SIZE = 4;
	defparam lut_1221.mask = 16'h1508;

	lut_sub lut_1223 ({sk[311], i_7_, i_32_, i_33_}, n_n861);
	defparam lut_1223.LUT_SIZE = 4;
	defparam lut_1223.mask = 16'h1540;

	lut_sub lut_1225 ({sk[312], i_39_, i_38_, i_37_}, n_n795);
	defparam lut_1225.LUT_SIZE = 4;
	defparam lut_1225.mask = 16'h1504;

	lut_sub lut_1227 ({sk[313], i_40_, i_39_, i_38_, i_37_}, x330x);
	defparam lut_1227.LUT_SIZE = 5;
	defparam lut_1227.mask = 32'h00ff0004;

	lut_sub lut_1229 ({sk[314], i_7_, i_32_, i_34_, i_33_, i_36_, i_35_}, x358x);
	defparam lut_1229.LUT_SIZE = 7;
	defparam lut_1229.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_1231 ({sk[315], i_34_, i_36_, i_35_}, n_n991);
	defparam lut_1231.LUT_SIZE = 4;
	defparam lut_1231.mask = 16'h1520;

	lut_sub lut_1233 ({sk[316], i_36_, i_35_}, x326x);
	defparam lut_1233.LUT_SIZE = 3;
	defparam lut_1233.mask = 8'h32;

	lut_sub lut_1235 ({sk[317], i_40_, i_7_, i_32_, i_34_, i_33_, x326x}, x435x);
	defparam lut_1235.LUT_SIZE = 7;
	defparam lut_1235.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_1237 ({sk[318], i_40_, i_34_, i_36_, i_35_}, x94x);
	defparam lut_1237.LUT_SIZE = 5;
	defparam lut_1237.mask = 32'h00ff0040;

	lut_sub lut_1239 ({sk[319], i_40_, i_7_, i_32_, i_33_, n_n979}, x528x);
	defparam lut_1239.LUT_SIZE = 6;
	defparam lut_1239.mask = 64'h55ffffff00001000;

	lut_sub lut_1241 ({sk[320], i_36_, i_38_, i_37_}, n_n1061);
	defparam lut_1241.LUT_SIZE = 4;
	defparam lut_1241.mask = 16'h1502;

	lut_sub lut_1243 ({sk[321], i_32_, i_34_, i_33_, i_35_}, x50x);
	defparam lut_1243.LUT_SIZE = 5;
	defparam lut_1243.mask = 32'h00ff1000;

	lut_sub lut_1245 ({sk[322], i_36_, i_38_, i_37_}, n_n582);
	defparam lut_1245.LUT_SIZE = 4;
	defparam lut_1245.mask = 16'h1510;

	lut_sub lut_1247 ({sk[323], i_40_, i_39_, i_38_, i_37_}, x400x);
	defparam lut_1247.LUT_SIZE = 5;
	defparam lut_1247.mask = 32'h00ff0002;

	lut_sub lut_1249 ({sk[324], i_32_, i_31_, i_33_, x109x, n_n1047, x400x}, n_n1373);
	defparam lut_1249.LUT_SIZE = 7;
	defparam lut_1249.mask = 128'h77777f7f77777f7f0001000000000000;

	lut_sub lut_1251 ({sk[325], i_30_, i_28_, i_29_}, x668x);
	defparam lut_1251.LUT_SIZE = 4;
	defparam lut_1251.mask = 16'h15db;

	lut_sub lut_1256 ({sk[326], i_40_, i_5_, i_39_, i_13_, i_15_}, x6783x);
	defparam lut_1256.LUT_SIZE = 6;
	defparam lut_1256.mask = 64'h55ffffff00008000;

	lut_sub lut_1258 ({sk[327], i_5_, x51x, x366x, n_n1048, x668x, x6783x}, x6784x);
	defparam lut_1258.LUT_SIZE = 7;
	defparam lut_1258.mask = 128'h77777f7f77777f7f0003555700005555;

	lut_sub lut_1261 ({sk[328], i_32_, i_31_, i_34_, i_33_, i_36_, i_35_}, x93x);
	defparam lut_1261.LUT_SIZE = 7;
	defparam lut_1261.mask = 128'h77777f7f77777f7f0800000000000000;

	lut_sub lut_1263 ({sk[329], i_39_, i_38_, i_37_}, n_n1001);
	defparam lut_1263.LUT_SIZE = 4;
	defparam lut_1263.mask = 16'h1502;

	lut_sub lut_1265 ({sk[330], i_3_, i_4_, i_1_, i_2_, x46x, n_n998}, n_n902);
	defparam lut_1265.LUT_SIZE = 7;
	defparam lut_1265.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_1267 ({sk[331], i_40_, i_5_, i_39_, i_38_}, x458x);
	defparam lut_1267.LUT_SIZE = 5;
	defparam lut_1267.mask = 32'h00ff0040;

	lut_sub lut_1269 ({sk[332], i_30_, i_28_, i_29_}, x669x);
	defparam lut_1269.LUT_SIZE = 4;
	defparam lut_1269.mask = 16'h155b;

	lut_sub lut_1273 ({sk[333], x6784x, x93x, n_n1001, n_n902, x458x, x669x}, n_n1164);
	defparam lut_1273.LUT_SIZE = 7;
	defparam lut_1273.mask = 128'h77777f7f77777f7f000f111fffffffff;

	lut_sub lut_1277 ({sk[334], i_40_, i_39_, i_21_, i_38_, x52x, x380x}, x1844x);
	defparam lut_1277.LUT_SIZE = 7;
	defparam lut_1277.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_1279 ({sk[335], n_n979, n_n945, n_n949, n_n947, n_n528, x399x}, x1846x);
	defparam lut_1279.LUT_SIZE = 7;
	defparam lut_1279.mask = 128'h77777f7f77777f7f0000000011111333;

	lut_sub lut_1283 ({sk[336], i_12_, i_11_, i_31_, x46x, n_n775, x407x}, x6793x);
	defparam lut_1283.LUT_SIZE = 7;
	defparam lut_1283.mask = 128'h77777f7f77777f7f0000010001000000;

	lut_sub lut_1286 ({sk[337], i_28_, i_29_, x93x, n_n902, x342x, x458x}, x6794x);
	defparam lut_1286.LUT_SIZE = 7;
	defparam lut_1286.mask = 128'h77777f7f77777f7f0357030303030303;

	lut_sub lut_1289 ({sk[338], i_21_, i_15_}, x48x);
	defparam lut_1289.LUT_SIZE = 3;
	defparam lut_1289.mask = 8'h34;

	lut_sub lut_1291 ({sk[339], i_5_, i_12_, i_11_, i_18_, i_15_}, x380x);
	defparam lut_1291.LUT_SIZE = 6;
	defparam lut_1291.mask = 64'h55ffffff01110000;

	lut_sub lut_1294 ({sk[340], i_9_, i_5_, i_12_, i_21_, i_15_, x380x}, x72x);
	defparam lut_1294.LUT_SIZE = 7;
	defparam lut_1294.mask = 128'h77777f7f77777f7f5050505050705050;

	lut_sub lut_1297 ({sk[341], i_40_, i_39_, i_32_, i_34_, i_33_}, x6797x);
	defparam lut_1297.LUT_SIZE = 6;
	defparam lut_1297.mask = 64'h55ffffff00004000;

	lut_sub lut_1299 ({sk[342], i_16_, i_32_, i_31_, i_33_, n_n1055, n_n1047}, x416x);
	defparam lut_1299.LUT_SIZE = 7;
	defparam lut_1299.mask = 128'h77777f7f77777f7f0000000001000000;

	lut_sub lut_1301 ({sk[343], i_12_, i_15_}, x78x);
	defparam lut_1301.LUT_SIZE = 3;
	defparam lut_1301.mask = 8'h31;

	lut_sub lut_1303 ({sk[344], i_17_, i_16_, n_n775, n_n1048, x98x, x522x}, x1835x);
	defparam lut_1303.LUT_SIZE = 7;
	defparam lut_1303.mask = 128'h77777f7f77777f7f0000000300070007;

	lut_sub lut_1307 ({sk[345], i_11_, x317x, n_n1372, x416x, x78x, x1835x}, x247x);
	defparam lut_1307.LUT_SIZE = 7;
	defparam lut_1307.mask = 128'h77777f7f77777f7f55ff57ff55ff55ff;

	lut_sub lut_1311 ({sk[346], i_36_, i_35_, i_37_}, n_n970);
	defparam lut_1311.LUT_SIZE = 4;
	defparam lut_1311.mask = 16'h1504;

	lut_sub lut_1313 ({sk[347], i_32_, i_34_, i_33_, i_36_, i_35_, i_37_}, x389x);
	defparam lut_1313.LUT_SIZE = 7;
	defparam lut_1313.mask = 128'h77777f7f77777f7f0004000000000000;

	lut_sub lut_1315 ({sk[348], i_39_, i_36_, i_35_, i_38_, i_37_, n_n1074}, x432x);
	defparam lut_1315.LUT_SIZE = 7;
	defparam lut_1315.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_1317 ({sk[349], i_23_, i_24_, i_22_}, n_n411);
	defparam lut_1317.LUT_SIZE = 4;
	defparam lut_1317.mask = 16'h1501;

	lut_sub lut_1319 ({sk[350], i_23_, i_24_, i_22_, i_19_}, x491x);
	defparam lut_1319.LUT_SIZE = 5;
	defparam lut_1319.mask = 32'h00ff0001;

	lut_sub lut_1321 ({sk[351], i_9_, i_5_, i_12_, i_11_, i_18_, i_19_}, x57x);
	defparam lut_1321.LUT_SIZE = 7;
	defparam lut_1321.mask = 128'h77777f7f77777f7f0000000007370000;

	lut_sub lut_1325 ({sk[352], i_39_, i_38_, x90x, n_n411, x57x}, x1831x);
	defparam lut_1325.LUT_SIZE = 6;
	defparam lut_1325.mask = 64'h55ffffff01000000;

	lut_sub lut_1327 ({sk[353], i_40_, i_38_}, n_n880);
	defparam lut_1327.LUT_SIZE = 3;
	defparam lut_1327.mask = 8'h32;

	lut_sub lut_1329 ({sk[354], i_3_, i_4_, i_1_, x314x, n_n926, n_n833}, x6818x);
	defparam lut_1329.LUT_SIZE = 7;
	defparam lut_1329.mask = 128'h77777f7f77777f7f0005050507070707;

	lut_sub lut_1334 ({sk[355], x88x, n_n991, x328x, x6811x, x325x, n_n997}, x6813x);
	defparam lut_1334.LUT_SIZE = 7;
	defparam lut_1334.mask = 128'h77777f7f77777f7f003300330f3f5f7f;

	lut_sub lut_1338 ({sk[356], i_40_, i_39_, i_38_}, n_n978);
	defparam lut_1338.LUT_SIZE = 4;
	defparam lut_1338.mask = 16'h1508;

	lut_sub lut_1340 ({sk[357], i_40_, i_39_, i_38_}, n_n883);
	defparam lut_1340.LUT_SIZE = 4;
	defparam lut_1340.mask = 16'h1504;

	lut_sub lut_1342 ({sk[358], i_36_, i_35_}, n_n964);
	defparam lut_1342.LUT_SIZE = 3;
	defparam lut_1342.mask = 8'h38;

	lut_sub lut_1344 ({sk[359], i_34_, i_36_, i_35_}, n_n998);
	defparam lut_1344.LUT_SIZE = 4;
	defparam lut_1344.mask = 16'h1508;

	lut_sub lut_1346 ({sk[360], i_7_, i_5_}, x47x);
	defparam lut_1346.LUT_SIZE = 3;
	defparam lut_1346.mask = 8'h38;

	lut_sub lut_1348 ({sk[361], i_7_, i_5_, i_13_}, n_n330);
	defparam lut_1348.LUT_SIZE = 4;
	defparam lut_1348.mask = 16'h1540;

	lut_sub lut_1350 ({sk[362], i_40_, i_39_, i_38_}, n_n969);
	defparam lut_1350.LUT_SIZE = 4;
	defparam lut_1350.mask = 16'h1580;

	lut_sub lut_1352 ({sk[363], i_9_, i_7_, i_5_, i_39_, i_38_, i_37_}, x6819x);
	defparam lut_1352.LUT_SIZE = 7;
	defparam lut_1352.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_1354 ({sk[364], i_15_, i_32_, i_33_}, n_n158);
	defparam lut_1354.LUT_SIZE = 4;
	defparam lut_1354.mask = 16'h1504;

	lut_sub lut_1356 ({sk[365], i_40_, i_9_, i_7_, i_5_, i_39_, i_38_}, x6820x);
	defparam lut_1356.LUT_SIZE = 7;
	defparam lut_1356.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_1358 ({sk[366], i_7_, i_32_, i_34_, i_33_, n_n964, n_n710}, n_n287);
	defparam lut_1358.LUT_SIZE = 7;
	defparam lut_1358.mask = 128'h77777f7f77777f7f0001000000000000;

	lut_sub lut_1360 ({sk[367], i_7_, i_3_, i_4_, i_0_, n_n1074, x95x}, x1805x);
	defparam lut_1360.LUT_SIZE = 7;
	defparam lut_1360.mask = 128'h77777f7f77777f7f0100010100000000;

	lut_sub lut_1363 ({sk[368], i_25_, i_26_, n_n864, n_n1011, x79x, x182x}, x6829x);
	defparam lut_1363.LUT_SIZE = 7;
	defparam lut_1363.mask = 128'h77777f7f77777f7f5557555555555555;

	lut_sub lut_1366 ({sk[369], x358x, n_n330, x100x, n_n710, n_n993, x6826x}, x6830x);
	defparam lut_1366.LUT_SIZE = 7;
	defparam lut_1366.mask = 128'h77777f7f77777f7f00001111000f111f;

	lut_sub lut_1369 ({sk[370], n_n785, x87x, x6852x, x1780x, x1781x, x8543x}, n_n1093);
	defparam lut_1369.LUT_SIZE = 7;
	defparam lut_1369.mask = 128'h77777f7f77777f7fbfbfbfbfbfbfbfff;

	lut_sub lut_1374 ({sk[371], n_n2793, x300x, x236x, x1765x, x1766x, x6868x}, n_n1091);
	defparam lut_1374.LUT_SIZE = 7;
	defparam lut_1374.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_1381 ({sk[372], x93x, x367x, x6859x, n_n1118, x6861x, x6877x}, x6879x);
	defparam lut_1381.LUT_SIZE = 7;
	defparam lut_1381.mask = 128'h77777f7f77777f7f7f7f7f7f7f7f7fff;

	lut_sub lut_1386 ({sk[373], i_39_, i_36_, x316x, n_n760, n_n764, x6875x}, x6878x);
	defparam lut_1386.LUT_SIZE = 7;
	defparam lut_1386.mask = 128'h77777f7f77777f7f55555555557f5555;

	lut_sub lut_1390 ({sk[374], x386x, x132x, x1717x, x6909x, x6910x}, x6913x);
	defparam lut_1390.LUT_SIZE = 6;
	defparam lut_1390.mask = 64'h55ffffff7f7f7fff;

	lut_sub lut_1395 ({sk[375], i_0_, i_36_, i_38_, i_37_}, x6920x);
	defparam lut_1395.LUT_SIZE = 5;
	defparam lut_1395.mask = 32'h00ff0010;

	lut_sub lut_1397 ({sk[376], i_7_, i_5_, i_11_}, n_n853);
	defparam lut_1397.LUT_SIZE = 4;
	defparam lut_1397.mask = 16'h1540;

	lut_sub lut_1399 ({sk[377], i_36_, i_35_, i_37_}, n_n968);
	defparam lut_1399.LUT_SIZE = 4;
	defparam lut_1399.mask = 16'h1520;

	lut_sub lut_1401 ({sk[378], i_40_, i_36_, i_35_, i_38_, i_37_}, x95x);
	defparam lut_1401.LUT_SIZE = 6;
	defparam lut_1401.mask = 64'h55ffffff00040000;

	lut_sub lut_1403 ({sk[379], i_7_, i_5_, i_13_, i_15_, x46x, n_n979}, x385x);
	defparam lut_1403.LUT_SIZE = 7;
	defparam lut_1403.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_1405 ({sk[380], i_40_, i_39_, i_38_, i_37_}, n_n469);
	defparam lut_1405.LUT_SIZE = 5;
	defparam lut_1405.mask = 32'h00ff0200;

	lut_sub lut_1407 ({sk[381], i_30_, i_7_, i_5_, i_28_, i_29_}, x6834x);
	defparam lut_1407.LUT_SIZE = 6;
	defparam lut_1407.mask = 64'h55ffffff00004000;

	lut_sub lut_1409 ({sk[382], i_40_, i_39_, i_38_}, n_n799);
	defparam lut_1409.LUT_SIZE = 4;
	defparam lut_1409.mask = 16'h1520;

	lut_sub lut_1411 ({sk[383], i_30_, i_7_, i_5_, i_28_, i_29_}, x6862x);
	defparam lut_1411.LUT_SIZE = 6;
	defparam lut_1411.mask = 64'h55ffffff20000000;

	lut_sub lut_1413 ({sk[384], i_39_, i_34_, i_36_, i_35_, i_38_, i_37_}, x6811x);
	defparam lut_1413.LUT_SIZE = 7;
	defparam lut_1413.mask = 128'h77777f7f77777f7f0000000000040000;

	lut_sub lut_1415 ({sk[385], i_32_, i_31_, i_34_, i_33_}, x76x);
	defparam lut_1415.LUT_SIZE = 5;
	defparam lut_1415.mask = 32'h00ff4000;

	lut_sub lut_1417 ({sk[386], i_24_, i_32_, i_33_}, n_n945);
	defparam lut_1417.LUT_SIZE = 4;
	defparam lut_1417.mask = 16'h1504;

	lut_sub lut_1419 ({sk[387], i_24_, i_22_, i_32_, i_33_, n_n979}, x52x);
	defparam lut_1419.LUT_SIZE = 6;
	defparam lut_1419.mask = 64'h55ffffff00000010;

	lut_sub lut_1421 ({sk[388], i_7_, i_5_, i_12_, i_21_, i_15_}, x329x);
	defparam lut_1421.LUT_SIZE = 6;
	defparam lut_1421.mask = 64'h55ffffff04000000;

	lut_sub lut_1423 ({sk[389], i_40_, i_39_, i_38_, i_37_}, x304x);
	defparam lut_1423.LUT_SIZE = 5;
	defparam lut_1423.mask = 32'h00ff8000;

	lut_sub lut_1425 ({sk[390], i_39_, i_34_, i_36_, i_35_, i_38_, i_37_}, x6939x);
	defparam lut_1425.LUT_SIZE = 7;
	defparam lut_1425.mask = 128'h77777f7f77777f7f0000008000000000;

	lut_sub lut_1427 ({sk[391], i_10_, i_27_, i_36_, i_35_, i_37_}, x6895x);
	defparam lut_1427.LUT_SIZE = 6;
	defparam lut_1427.mask = 64'h55ffffff00000008;

	lut_sub lut_1429 ({sk[392], i_23_, i_21_, i_15_, x90x, n_n978, n_n850}, x1691x);
	defparam lut_1429.LUT_SIZE = 7;
	defparam lut_1429.mask = 128'h77777f7f77777f7f0001000000000000;

	lut_sub lut_1431 ({sk[393], i_39_, i_38_, i_37_, n_n1047, x87x, x6852x}, x1692x);
	defparam lut_1431.LUT_SIZE = 7;
	defparam lut_1431.mask = 128'h77777f7f77777f7f0001000000000000;

	lut_sub lut_1433 ({sk[394], i_31_, n_n1074, n_n1012, n_n799, x6834x, x6862x}, x6940x);
	defparam lut_1433.LUT_SIZE = 7;
	defparam lut_1433.mask = 128'h77777f7f77777f7f0000000700000000;

	lut_sub lut_1436 ({sk[395], i_32_, n_n1008, n_n1052, x365x, n_n2456, n_n1023}, x6941x);
	defparam lut_1436.LUT_SIZE = 7;
	defparam lut_1436.mask = 128'h77777f7f77777f7f3333333733333333;

	lut_sub lut_1439 ({sk[396], n_n880, n_n960, n_n1047, n_n2793, x368x, x6850x}, x6942x);
	defparam lut_1439.LUT_SIZE = 7;
	defparam lut_1439.mask = 128'h77777f7f77777f7f0f0f0f1f0f1f0f1f;

	lut_sub lut_1443 ({sk[397], i_40_, i_39_, i_36_, i_38_, n_n837}, x1682x);
	defparam lut_1443.LUT_SIZE = 6;
	defparam lut_1443.mask = 64'h55ffffff00004000;

	lut_sub lut_1445 ({sk[398], i_39_, i_36_, i_38_, i_37_, n_n760, n_n834}, x6946x);
	defparam lut_1445.LUT_SIZE = 7;
	defparam lut_1445.mask = 128'h77777f7f77777f7f5000000000300000;

	lut_sub lut_1448 ({sk[399], i_39_, i_38_, n_n1047, x68x, x367x, x6858x}, n_n1118);
	defparam lut_1448.LUT_SIZE = 7;
	defparam lut_1448.mask = 128'h77777f7f77777f7f0001000100010011;

	lut_sub lut_1451 ({sk[400], i_22_, i_32_, x82x, x359x, x101x, n_n1023}, x1675x);
	defparam lut_1451.LUT_SIZE = 7;
	defparam lut_1451.mask = 128'h77777f7f77777f7f0015000000000000;

	lut_sub lut_1454 ({sk[401], i_40_, i_39_, n_n985, x365x, n_n1980, x80x}, x6950x);
	defparam lut_1454.LUT_SIZE = 7;
	defparam lut_1454.mask = 128'h77777f7f77777f7f3333333333333337;

	lut_sub lut_1457 ({sk[402], i_23_, i_32_, x82x, x323x, x365x, n_n1023}, x6951x);
	defparam lut_1457.LUT_SIZE = 7;
	defparam lut_1457.mask = 128'h77777f7f77777f7f0105000001010000;

	lut_sub lut_1460 ({sk[403], i_22_, i_32_, i_34_, i_33_, i_35_, x82x}, n_n764);
	defparam lut_1460.LUT_SIZE = 7;
	defparam lut_1460.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_1462 ({sk[404], i_24_, i_32_, x82x, x54x, n_n1023}, x240x);
	defparam lut_1462.LUT_SIZE = 6;
	defparam lut_1462.mask = 64'h55ffffff01000000;

	lut_sub lut_1464 ({sk[405], n_n1935, n_n1936, x6958x, x6956x, x6957x}, x8542x);
	defparam lut_1464.LUT_SIZE = 6;
	defparam lut_1464.mask = 64'h55ffffff80000000;

	lut_sub lut_1466 ({sk[406], i_24_, i_32_, i_34_, i_33_, i_35_, x87x}, n_n834);
	defparam lut_1466.LUT_SIZE = 7;
	defparam lut_1466.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_1468 ({sk[407], i_39_, i_36_, i_38_}, n_n836);
	defparam lut_1468.LUT_SIZE = 4;
	defparam lut_1468.mask = 16'h1580;

	lut_sub lut_1470 ({sk[408], i_40_, n_n861, x6811x, n_n833, n_n834, n_n836}, x173x);
	defparam lut_1470.LUT_SIZE = 7;
	defparam lut_1470.mask = 128'h77777f7f77777f7f030303ff13131313;

	lut_sub lut_1474 ({sk[409], i_9_, i_7_, i_5_}, n_n793);
	defparam lut_1474.LUT_SIZE = 4;
	defparam lut_1474.mask = 16'h1580;

	lut_sub lut_1476 ({sk[410], i_40_, i_39_, i_38_, i_37_, x93x, n_n793}, x181x);
	defparam lut_1476.LUT_SIZE = 7;
	defparam lut_1476.mask = 128'h77777f7f77777f7f0000001100000001;

	lut_sub lut_1479 ({sk[411], i_7_, i_5_, i_11_, i_15_}, x82x);
	defparam lut_1479.LUT_SIZE = 5;
	defparam lut_1479.mask = 32'h00ff1000;

	lut_sub lut_1481 ({sk[412], i_7_, i_5_, i_12_, i_15_}, x87x);
	defparam lut_1481.LUT_SIZE = 5;
	defparam lut_1481.mask = 32'h00ff1000;

	lut_sub lut_1483 ({sk[413], i_17_, i_16_}, x37x);
	defparam lut_1483.LUT_SIZE = 3;
	defparam lut_1483.mask = 8'h37;

	lut_sub lut_1486 ({sk[414], i_40_, x368x, x367x, x6976x, x6977x, x1657x}, x1653x);
	defparam lut_1486.LUT_SIZE = 7;
	defparam lut_1486.mask = 128'h77777f7f77777f7f0000000001030303;

	lut_sub lut_1490 ({sk[415], i_18_, n_n1055, x94x, x368x, n_n791, x367x}, x1652x);
	defparam lut_1490.LUT_SIZE = 7;
	defparam lut_1490.mask = 128'h77777f7f77777f7f0000001300000000;

	lut_sub lut_1493 ({sk[416], i_16_, i_31_, x46x, x368x, x64x, x367x}, x1661x);
	defparam lut_1493.LUT_SIZE = 7;
	defparam lut_1493.mask = 128'h77777f7f77777f7f0013000000000000;

	lut_sub lut_1496 ({sk[417], i_17_, i_31_, x46x, n_n775, x368x, x367x}, x6970x);
	defparam lut_1496.LUT_SIZE = 7;
	defparam lut_1496.mask = 128'h77777f7f77777f7f0007000000000000;

	lut_sub lut_1499 ({sk[418], n_n979, n_n1001, n_n775, x367x, n_n773, x6968x}, x6971x);
	defparam lut_1499.LUT_SIZE = 7;
	defparam lut_1499.mask = 128'h77777f7f77777f7f0033003300330537;

	lut_sub lut_1502 ({sk[419], i_23_, n_n979, n_n1001, x365x, n_n857, n_n790}, x8541x);
	defparam lut_1502.LUT_SIZE = 7;
	defparam lut_1502.mask = 128'h77777f7f77777f7ffcfcfca8ffffffaa;

	lut_sub lut_1512 ({sk[420], i_7_, i_5_, i_0_}, n_n685);
	defparam lut_1512.LUT_SIZE = 4;
	defparam lut_1512.mask = 16'h1520;

	lut_sub lut_1514 ({sk[421], i_7_, i_39_, i_36_, i_38_, i_37_, x80x}, x438x);
	defparam lut_1514.LUT_SIZE = 7;
	defparam lut_1514.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_1516 ({sk[422], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x431x);
	defparam lut_1516.LUT_SIZE = 7;
	defparam lut_1516.mask = 128'h77777f7f77777f7f0000000000100000;

	lut_sub lut_1518 ({sk[423], i_7_, i_1_, i_0_, i_32_, i_34_, i_33_}, x541x);
	defparam lut_1518.LUT_SIZE = 7;
	defparam lut_1518.mask = 128'h77777f7f77777f7f0000004000000000;

	lut_sub lut_1520 ({sk[424], i_7_, i_0_, i_32_, i_34_, i_33_}, x350x);
	defparam lut_1520.LUT_SIZE = 6;
	defparam lut_1520.mask = 64'h55ffffff00400000;

	lut_sub lut_1522 ({sk[425], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x362x);
	defparam lut_1522.LUT_SIZE = 7;
	defparam lut_1522.mask = 128'h77777f7f77777f7f0000000000000020;

	lut_sub lut_1524 ({sk[426], i_40_, i_39_, i_36_, x316x, x7006x, n_n1023}, x341x);
	defparam lut_1524.LUT_SIZE = 7;
	defparam lut_1524.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_1526 ({sk[427], i_7_, i_5_, i_12_, i_11_, i_18_}, x412x);
	defparam lut_1526.LUT_SIZE = 6;
	defparam lut_1526.mask = 64'h55ffffff15000000;

	lut_sub lut_1529 ({sk[428], i_17_, i_32_, i_31_, i_34_, i_33_, i_35_}, x425x);
	defparam lut_1529.LUT_SIZE = 7;
	defparam lut_1529.mask = 128'h77777f7f77777f7f0000000020000000;

	lut_sub lut_1531 ({sk[429], i_17_, i_32_, i_31_}, n_n933);
	defparam lut_1531.LUT_SIZE = 4;
	defparam lut_1531.mask = 16'h1508;

	lut_sub lut_1533 ({sk[430], i_32_, i_33_, i_35_}, n_n874);
	defparam lut_1533.LUT_SIZE = 4;
	defparam lut_1533.mask = 16'h1520;

	lut_sub lut_1535 ({sk[431], i_32_, i_31_, i_33_, i_35_}, x422x);
	defparam lut_1535.LUT_SIZE = 5;
	defparam lut_1535.mask = 32'h00ff2000;

	lut_sub lut_1537 ({sk[432], i_40_, i_39_, i_36_, i_38_}, n_n462);
	defparam lut_1537.LUT_SIZE = 5;
	defparam lut_1537.mask = 32'h00ff0040;

	lut_sub lut_1539 ({sk[433], i_30_, i_7_, i_5_, i_28_, i_29_}, x7019x);
	defparam lut_1539.LUT_SIZE = 6;
	defparam lut_1539.mask = 64'h55ffffff80000000;

	lut_sub lut_1541 ({sk[434], i_7_, i_5_, i_11_}, n_n527);
	defparam lut_1541.LUT_SIZE = 4;
	defparam lut_1541.mask = 16'h1580;

	lut_sub lut_1543 ({sk[435], i_16_, i_32_, i_31_, i_34_, i_33_, i_35_}, x388x);
	defparam lut_1543.LUT_SIZE = 7;
	defparam lut_1543.mask = 128'h77777f7f77777f7f0000000020000000;

	lut_sub lut_1545 ({sk[436], i_9_, i_7_, i_5_, i_12_, i_11_, i_15_}, x7015x);
	defparam lut_1545.LUT_SIZE = 7;
	defparam lut_1545.mask = 128'h77777f7f77777f7f0000000014000000;

	lut_sub lut_1548 ({sk[437], i_34_, i_33_, i_35_}, n_n1023);
	defparam lut_1548.LUT_SIZE = 4;
	defparam lut_1548.mask = 16'h1510;

	lut_sub lut_1550 ({sk[438], i_21_, i_15_, i_32_, n_n850, n_n1023}, n_n761);
	defparam lut_1550.LUT_SIZE = 6;
	defparam lut_1550.mask = 64'h55ffffff00100000;

	lut_sub lut_1552 ({sk[439], i_22_, i_32_, i_34_, i_33_, i_35_, x87x}, n_n760);
	defparam lut_1552.LUT_SIZE = 7;
	defparam lut_1552.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_1554 ({sk[440], i_40_, i_39_, i_36_, x81x, x329x, x80x}, n_n1928);
	defparam lut_1554.LUT_SIZE = 7;
	defparam lut_1554.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_1556 ({sk[441], i_40_, i_39_, i_22_, n_n985, x80x, x87x}, n_n1983);
	defparam lut_1556.LUT_SIZE = 7;
	defparam lut_1556.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_1558 ({sk[442], i_40_, i_39_, i_23_, i_36_, i_38_, i_37_}, x6955x);
	defparam lut_1558.LUT_SIZE = 7;
	defparam lut_1558.mask = 128'h77777f7f77777f7f0000200000000000;

	lut_sub lut_1560 ({sk[443], i_40_, i_39_, i_36_, i_38_, i_37_}, x359x);
	defparam lut_1560.LUT_SIZE = 6;
	defparam lut_1560.mask = 64'h55ffffff00004000;

	lut_sub lut_1562 ({sk[444], i_40_, i_39_, i_36_, i_38_, i_37_}, x101x);
	defparam lut_1562.LUT_SIZE = 6;
	defparam lut_1562.mask = 64'h55ffffff80000000;

	lut_sub lut_1564 ({sk[445], i_17_, i_16_, n_n960, n_n1047, n_n1048, x367x}, x174x);
	defparam lut_1564.LUT_SIZE = 7;
	defparam lut_1564.mask = 128'h77777f7f77777f7f0001000100010000;

	lut_sub lut_1567 ({sk[446], x329x, x50x, n_n764, x359x, x101x, x174x}, x7028x);
	defparam lut_1567.LUT_SIZE = 7;
	defparam lut_1567.mask = 128'h77777f7f77777f7f557f557f557f777f;

	lut_sub lut_1572 ({sk[447], i_40_, i_39_, i_22_, n_n985, x82x, x80x}, n_n1980);
	defparam lut_1572.LUT_SIZE = 7;
	defparam lut_1572.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_1574 ({sk[448], i_40_, i_39_, i_38_, i_37_}, x68x);
	defparam lut_1574.LUT_SIZE = 5;
	defparam lut_1574.mask = 32'h00ff0ace;

	lut_sub lut_1577 ({sk[449], i_16_, i_34_, i_36_, i_35_, n_n1048, x367x}, x504x);
	defparam lut_1577.LUT_SIZE = 7;
	defparam lut_1577.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_1579 ({sk[450], i_23_, i_32_, x82x, x323x, n_n1023}, x157x);
	defparam lut_1579.LUT_SIZE = 6;
	defparam lut_1579.mask = 64'h55ffffff01000000;

	lut_sub lut_1581 ({sk[451], i_40_, i_39_, i_36_, x81x, x365x, x80x}, n_n1927);
	defparam lut_1581.LUT_SIZE = 7;
	defparam lut_1581.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_1583 ({sk[452], i_39_, i_34_, i_37_, n_n964, x368x, x6850x}, n_n2793);
	defparam lut_1583.LUT_SIZE = 7;
	defparam lut_1583.mask = 128'h77777f7f77777f7f0000000001000000;

	lut_sub lut_1585 ({sk[453], i_39_, i_17_, i_38_, n_n1047, n_n1048, x368x}, n_n2456);
	defparam lut_1585.LUT_SIZE = 7;
	defparam lut_1585.mask = 128'h77777f7f77777f7f0000000000010000;

	lut_sub lut_1587 ({sk[454], i_40_, i_39_, i_38_, n_n1047, x368x, x6850x}, x300x);
	defparam lut_1587.LUT_SIZE = 7;
	defparam lut_1587.mask = 128'h77777f7f77777f7f0000000101000101;

	lut_sub lut_1590 ({sk[455], n_n1008, x323x, n_n1052, n_n765, x1691x, x1692x}, x8539x);
	defparam lut_1590.LUT_SIZE = 7;
	defparam lut_1590.mask = 128'h77777f7f77777f7f8888808088808080;

	lut_sub lut_1594 ({sk[456], i_40_, i_39_, i_36_, i_38_, i_37_}, x323x);
	defparam lut_1594.LUT_SIZE = 6;
	defparam lut_1594.mask = 64'h55ffffff00200000;

	lut_sub lut_1596 ({sk[457], i_39_, i_38_, i_37_}, n_n975);
	defparam lut_1596.LUT_SIZE = 4;
	defparam lut_1596.mask = 16'h1580;

	lut_sub lut_1598 ({sk[458], i_1_, i_2_, i_0_}, n_n843);
	defparam lut_1598.LUT_SIZE = 4;
	defparam lut_1598.mask = 16'h1510;

	lut_sub lut_1600 ({sk[459], i_5_, i_32_, i_33_}, n_n980);
	defparam lut_1600.LUT_SIZE = 4;
	defparam lut_1600.mask = 16'h1504;

	lut_sub lut_1602 ({sk[460], i_5_, i_0_, i_32_}, n_n1006);
	defparam lut_1602.LUT_SIZE = 4;
	defparam lut_1602.mask = 16'h1508;

	lut_sub lut_1604 ({sk[461], i_15_, i_32_, i_31_}, n_n989);
	defparam lut_1604.LUT_SIZE = 4;
	defparam lut_1604.mask = 16'h1580;

	lut_sub lut_1606 ({sk[462], i_34_, i_33_}, x322x);
	defparam lut_1606.LUT_SIZE = 3;
	defparam lut_1606.mask = 8'h34;

	lut_sub lut_1608 ({sk[463], i_34_, i_33_, i_36_}, n_n983);
	defparam lut_1608.LUT_SIZE = 4;
	defparam lut_1608.mask = 16'h1520;

	lut_sub lut_1610 ({sk[464], i_39_, i_38_, i_37_}, x65x);
	defparam lut_1610.LUT_SIZE = 4;
	defparam lut_1610.mask = 16'h1582;

	lut_sub lut_1613 ({sk[465], i_7_, i_34_, i_33_, i_36_, n_n980, x65x}, x7048x);
	defparam lut_1613.LUT_SIZE = 7;
	defparam lut_1613.mask = 128'h77777f7f77777f7f1010000010ff00ff;

	lut_sub lut_1616 ({sk[466], i_36_, i_38_, i_37_, n_n1023, n_n1057}, x518x);
	defparam lut_1616.LUT_SIZE = 6;
	defparam lut_1616.mask = 64'h55ffffff00000001;

	lut_sub lut_1618 ({sk[467], i_12_, i_11_, x76x, x327x, x110x, x827x}, x1567x);
	defparam lut_1618.LUT_SIZE = 7;
	defparam lut_1618.mask = 128'h77777f7f77777f7f005d000c000c000c;

	lut_sub lut_1621 ({sk[468], i_35_, i_37_, n_n977, x41x, x452x, x1566x}, x7061x);
	defparam lut_1621.LUT_SIZE = 7;
	defparam lut_1621.mask = 128'h77777f7f77777f7f5557555555555555;

	lut_sub lut_1624 ({sk[469], i_9_, i_12_, x84x, x76x, x37x, x327x}, x1575x);
	defparam lut_1624.LUT_SIZE = 7;
	defparam lut_1624.mask = 128'h77777f7f77777f7f0000000001330101;

	lut_sub lut_1627 ({sk[470], i_40_, i_39_, x45x, n_n1067, x393x, x8548x}, x1557x);
	defparam lut_1627.LUT_SIZE = 7;
	defparam lut_1627.mask = 128'h77777f7f77777f7f030b030b030b000a;

	lut_sub lut_1631 ({sk[471], i_40_, i_36_, n_n1159, n_n1055, x322x, x472x}, x7069x);
	defparam lut_1631.LUT_SIZE = 7;
	defparam lut_1631.mask = 128'h77777f7f77777f7f00ff01ff00ff00ff;

	lut_sub lut_1634 ({sk[472], i_9_, i_14_, i_11_, x84x, x416x, x7051x}, x8538x);
	defparam lut_1634.LUT_SIZE = 7;
	defparam lut_1634.mask = 128'h77777f7f77777f7ffafafafac8c8c8fa;

	lut_sub lut_1641 ({sk[473], i_15_, i_32_, i_31_, i_34_, i_33_, i_35_}, x387x);
	defparam lut_1641.LUT_SIZE = 7;
	defparam lut_1641.mask = 128'h77777f7f77777f7f2000000000000000;

	lut_sub lut_1643 ({sk[474], i_40_, i_39_, i_36_, i_38_, i_37_}, x119x);
	defparam lut_1643.LUT_SIZE = 6;
	defparam lut_1643.mask = 64'h55ffffff008000a0;

	lut_sub lut_1646 ({sk[475], i_40_, i_6_, x819x}, x1538x);
	defparam lut_1646.LUT_SIZE = 4;
	defparam lut_1646.mask = 16'h1501;

	lut_sub lut_1648 ({sk[476], i_36_, n_n1006, x322x, x441x, x397x, x7078x}, x7084x);
	defparam lut_1648.LUT_SIZE = 7;
	defparam lut_1648.mask = 128'h77777f7f77777f7f111111111111111f;

	lut_sub lut_1651 ({sk[477], i_12_, i_11_, i_31_, n_n1074, x401x, x1539x}, x7085x);
	defparam lut_1651.LUT_SIZE = 7;
	defparam lut_1651.mask = 128'h77777f7f77777f7f5755555555555555;

	lut_sub lut_1654 ({sk[478], i_40_, i_39_, i_38_, i_37_}, x445x);
	defparam lut_1654.LUT_SIZE = 5;
	defparam lut_1654.mask = 32'h00ff2000;

	lut_sub lut_1656 ({sk[479], i_33_, i_36_, i_35_}, n_n976);
	defparam lut_1656.LUT_SIZE = 4;
	defparam lut_1656.mask = 16'h1508;

	lut_sub lut_1658 ({sk[480], i_40_, i_39_, i_38_, i_37_, n_n1066, n_n976}, x7090x);
	defparam lut_1658.LUT_SIZE = 7;
	defparam lut_1658.mask = 128'h77777f7f77777f7f5000503050000030;

	lut_sub lut_1662 ({sk[481], i_36_, i_37_}, x355x);
	defparam lut_1662.LUT_SIZE = 3;
	defparam lut_1662.mask = 8'h31;

	lut_sub lut_1664 ({sk[482], i_7_, i_34_}, x453x);
	defparam lut_1664.LUT_SIZE = 3;
	defparam lut_1664.mask = 8'h38;

	lut_sub lut_1666 ({sk[483], i_34_, i_35_, i_37_}, n_n715);
	defparam lut_1666.LUT_SIZE = 4;
	defparam lut_1666.mask = 16'h1510;

	lut_sub lut_1668 ({sk[484], i_40_, i_39_, i_38_, i_37_, n_n998, n_n715}, x7104x);
	defparam lut_1668.LUT_SIZE = 7;
	defparam lut_1668.mask = 128'h77777f7f77777f7f3000305530000000;

	lut_sub lut_1672 ({sk[485], i_32_, i_34_, i_36_, i_35_, n_n709, n_n1008}, x1510x);
	defparam lut_1672.LUT_SIZE = 7;
	defparam lut_1672.mask = 128'h77777f7f77777f7f000000000ffff010;

	lut_sub lut_1677 ({sk[486], i_36_, i_35_, i_37_}, n_n971);
	defparam lut_1677.LUT_SIZE = 4;
	defparam lut_1677.mask = 16'h1508;

	lut_sub lut_1679 ({sk[487], i_38_, i_37_}, x100x);
	defparam lut_1679.LUT_SIZE = 3;
	defparam lut_1679.mask = 8'h31;

	lut_sub lut_1681 ({sk[488], i_39_, i_38_}, n_n960);
	defparam lut_1681.LUT_SIZE = 3;
	defparam lut_1681.mask = 8'h31;

	lut_sub lut_1683 ({sk[489], i_39_, i_38_, i_37_}, n_n997);
	defparam lut_1683.LUT_SIZE = 4;
	defparam lut_1683.mask = 16'h1501;

	lut_sub lut_1685 ({sk[490], i_7_, i_12_, i_11_, i_32_, i_34_, i_33_}, x390x);
	defparam lut_1685.LUT_SIZE = 7;
	defparam lut_1685.mask = 128'h77777f7f77777f7f4000000000000000;

	lut_sub lut_1687 ({sk[491], i_40_, i_7_, i_32_, i_34_, i_33_, n_n964}, x510x);
	defparam lut_1687.LUT_SIZE = 7;
	defparam lut_1687.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_1689 ({sk[492], i_7_, i_32_, i_34_, i_33_}, x79x);
	defparam lut_1689.LUT_SIZE = 5;
	defparam lut_1689.mask = 32'h00ff4000;

	lut_sub lut_1691 ({sk[493], i_7_, i_3_, i_4_, n_n1074, n_n1067}, x526x);
	defparam lut_1691.LUT_SIZE = 6;
	defparam lut_1691.mask = 64'h55ffffff10000000;

	lut_sub lut_1693 ({sk[494], i_32_, i_34_, i_33_}, n_n966);
	defparam lut_1693.LUT_SIZE = 4;
	defparam lut_1693.mask = 16'h1510;

	lut_sub lut_1695 ({sk[495], i_36_, i_35_, i_38_}, n_n862);
	defparam lut_1695.LUT_SIZE = 4;
	defparam lut_1695.mask = 16'h1540;

	lut_sub lut_1697 ({sk[496], i_39_, i_38_}, x346x);
	defparam lut_1697.LUT_SIZE = 3;
	defparam lut_1697.mask = 8'h34;

	lut_sub lut_1699 ({sk[497], o_15_, n_n1064, n_n966, n_n862, x346x, x89x}, x122x);
	defparam lut_1699.LUT_SIZE = 7;
	defparam lut_1699.mask = 128'h77777f7f77777f7f1111111fffffffff;

	lut_sub lut_1703 ({sk[498], i_7_, i_34_, i_33_, i_36_, i_35_}, x49x);
	defparam lut_1703.LUT_SIZE = 6;
	defparam lut_1703.mask = 64'h55ffffff08000000;

	lut_sub lut_1705 ({sk[499], i_9_, i_12_, i_11_, i_16_, i_15_}, x8571x);
	defparam lut_1705.LUT_SIZE = 6;
	defparam lut_1705.mask = 64'h55fffffffefefaaa;

	lut_sub lut_1710 ({sk[500], i_7_, i_31_, i_34_, i_33_, i_36_, i_35_}, x354x);
	defparam lut_1710.LUT_SIZE = 7;
	defparam lut_1710.mask = 128'h77777f7f77777f7f0800000000000000;

	lut_sub lut_1712 ({sk[501], i_11_, i_15_}, x86x);
	defparam lut_1712.LUT_SIZE = 3;
	defparam lut_1712.mask = 8'h31;

	lut_sub lut_1714 ({sk[502], i_9_, i_16_, n_n973, n_n967, x86x, x78x}, x8566x);
	defparam lut_1714.LUT_SIZE = 7;
	defparam lut_1714.mask = 128'h77777f7f77777f7ffffffcccfaaaf888;

	lut_sub lut_1729 ({sk[503], i_9_, n_n973, n_n967, x354x, x86x, x8566x}, x7210x);
	defparam lut_1729.LUT_SIZE = 7;
	defparam lut_1729.mask = 128'h77777f7f77777f7f0a0a0a0a0a0b0b0b;

	lut_sub lut_1733 ({sk[504], i_7_, i_5_, i_0_, i_32_, i_34_, i_33_}, x428x);
	defparam lut_1733.LUT_SIZE = 7;
	defparam lut_1733.mask = 128'h77777f7f77777f7f0000400000000000;

	lut_sub lut_1735 ({sk[505], i_40_, i_31_, n_n1066, x344x, x383x, x166x}, x1383x);
	defparam lut_1735.LUT_SIZE = 7;
	defparam lut_1735.mask = 128'h77777f7f77777f7f0002000000000000;

	lut_sub lut_1737 ({sk[506], i_7_, i_5_, i_32_, i_33_, i_36_, i_35_}, x7212x);
	defparam lut_1737.LUT_SIZE = 7;
	defparam lut_1737.mask = 128'h77777f7f77777f7f0000080000000000;

	lut_sub lut_1739 ({sk[507], i_7_, i_5_, i_32_}, n_n668);
	defparam lut_1739.LUT_SIZE = 4;
	defparam lut_1739.mask = 16'h1520;

	lut_sub lut_1741 ({sk[508], i_39_, i_36_, i_38_, i_37_, x322x, n_n668}, x251x);
	defparam lut_1741.LUT_SIZE = 7;
	defparam lut_1741.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_1743 ({sk[509], i_32_, i_34_, i_33_, i_36_, i_35_, i_37_}, x502x);
	defparam lut_1743.LUT_SIZE = 7;
	defparam lut_1743.mask = 128'h77777f7f77777f7f0001000000000000;

	lut_sub lut_1745 ({sk[510], i_36_, i_38_, i_37_}, n_n1052);
	defparam lut_1745.LUT_SIZE = 4;
	defparam lut_1745.mask = 16'h1580;

	lut_sub lut_1747 ({sk[511], i_32_, i_33_, i_36_, i_35_, n_n709, n_n685}, x392x);
	defparam lut_1747.LUT_SIZE = 7;
	defparam lut_1747.mask = 128'h77777f7f77777f7f0000100000000000;

	lut_sub lut_1749 ({sk[512], i_7_, i_5_, i_34_, i_33_, i_36_, i_35_}, x405x);
	defparam lut_1749.LUT_SIZE = 7;
	defparam lut_1749.mask = 128'h77777f7f77777f7f0000080000000000;

	lut_sub lut_1751 ({sk[513], i_40_, i_39_, i_37_}, n_n528);
	defparam lut_1751.LUT_SIZE = 4;
	defparam lut_1751.mask = 16'h1508;

	lut_sub lut_1753 ({sk[514], i_35_, n_n1014, n_n1074, n_n985, n_n975, n_n528}, x1364x);
	defparam lut_1753.LUT_SIZE = 7;
	defparam lut_1753.mask = 128'h77777f7f77777f7f000f0000007f0077;

	lut_sub lut_1757 ({sk[515], i_34_, i_35_}, x490x);
	defparam lut_1757.LUT_SIZE = 3;
	defparam lut_1757.mask = 8'h38;

	lut_sub lut_1759 ({sk[516], i_15_, i_32_, i_33_}, n_n700);
	defparam lut_1759.LUT_SIZE = 4;
	defparam lut_1759.mask = 16'h1540;

	lut_sub lut_1761 ({sk[517], n_n1008, n_n874, n_n1006, x322x, x100x, n_n693}, x7235x);
	defparam lut_1761.LUT_SIZE = 7;
	defparam lut_1761.mask = 128'h77777f7f77777f7f0003000300035557;

	lut_sub lut_1764 ({sk[518], i_9_, i_16_}, x404x);
	defparam lut_1764.LUT_SIZE = 3;
	defparam lut_1764.mask = 8'h38;

	lut_sub lut_1766 ({sk[519], i_12_, i_11_}, x61x);
	defparam lut_1766.LUT_SIZE = 3;
	defparam lut_1766.mask = 8'h37;

	lut_sub lut_1769 ({sk[520], i_32_, i_33_, i_36_, i_35_}, x421x);
	defparam lut_1769.LUT_SIZE = 5;
	defparam lut_1769.mask = 32'h00ff0800;

	lut_sub lut_1771 ({sk[521], x45x, x316x, n_n880, x404x, x61x, x421x}, x1349x);
	defparam lut_1771.LUT_SIZE = 7;
	defparam lut_1771.mask = 128'h77777f7f77777f7f0000454500cf45cf;

	lut_sub lut_1776 ({sk[522], i_32_, i_34_, i_33_, i_36_, i_35_}, x77x);
	defparam lut_1776.LUT_SIZE = 6;
	defparam lut_1776.mask = 64'h55ffffff00080000;

	lut_sub lut_1778 ({sk[523], i_3_, i_1_, i_2_, i_0_}, x464x);
	defparam lut_1778.LUT_SIZE = 5;
	defparam lut_1778.mask = 32'h00ff1000;

	lut_sub lut_1780 ({sk[524], n_n709, x45x, n_n1006, n_n976, x61x, n_n918}, x7259x);
	defparam lut_1780.LUT_SIZE = 7;
	defparam lut_1780.mask = 128'h77777f7f77777f7f00004444000f444f;

	lut_sub lut_1783 ({sk[525], i_32_, i_31_, i_34_, i_33_, i_36_, i_35_}, x339x);
	defparam lut_1783.LUT_SIZE = 7;
	defparam lut_1783.mask = 128'h77777f7f77777f7f0000080000000000;

	lut_sub lut_1785 ({sk[526], i_5_, i_32_, i_34_, i_33_, i_36_, i_35_}, x424x);
	defparam lut_1785.LUT_SIZE = 7;
	defparam lut_1785.mask = 128'h77777f7f77777f7f0000000008000000;

	lut_sub lut_1787 ({sk[527], i_31_, i_34_, i_33_, n_n860, x521x, x8528x}, x1308x);
	defparam lut_1787.LUT_SIZE = 7;
	defparam lut_1787.mask = 128'h77777f7f77777f7f00ab00aa00000000;

	lut_sub lut_1790 ({sk[528], i_40_, i_39_, n_n990, x328x, n_n888, x97x}, x7283x);
	defparam lut_1790.LUT_SIZE = 7;
	defparam lut_1790.mask = 128'h77777f7f77777f7f00000000111f000f;

	lut_sub lut_1793 ({sk[529], i_39_, i_37_, n_n861, n_n998, n_n710, x8527x}, x7284x);
	defparam lut_1793.LUT_SIZE = 7;
	defparam lut_1793.mask = 128'h77777f7f77777f7faaabaaaaaaaaaaaa;

	lut_sub lut_1796 ({sk[530], n_n883, n_n1047, n_n287, n_n799, x102x, x488x}, x7299x);
	defparam lut_1796.LUT_SIZE = 7;
	defparam lut_1796.mask = 128'h77777f7f77777f7f000f000f000f111f;

	lut_sub lut_1799 ({sk[531], i_40_, i_36_, i_38_, n_n515, x398x}, x8526x);
	defparam lut_1799.LUT_SIZE = 6;
	defparam lut_1799.mask = 64'h55fffffff8fafafa;

	lut_sub lut_1804 ({sk[532], n_n795, n_n1047, n_n535, n_n688, x488x, x765x}, x764x);
	defparam lut_1804.LUT_SIZE = 7;
	defparam lut_1804.mask = 128'h77777f7f77777f7f000f000f000f111f;

	lut_sub lut_1807 ({sk[533], i_24_, i_32_, n_n528, n_n525, n_n1023, x486x}, x1284x);
	defparam lut_1807.LUT_SIZE = 7;
	defparam lut_1807.mask = 128'h77777f7f77777f7f000f000f001f000f;

	lut_sub lut_1810 ({sk[534], i_16_, i_31_, x82x, n_n1066, n_n1052, x87x}, x1285x);
	defparam lut_1810.LUT_SIZE = 7;
	defparam lut_1810.mask = 128'h77777f7f77777f7f0000000001030000;

	lut_sub lut_1813 ({sk[535], i_31_, i_36_, n_n709, n_n1066, x7288x, x7289x}, x1293x);
	defparam lut_1813.LUT_SIZE = 7;
	defparam lut_1813.mask = 128'h77777f7f77777f7f0007000000000000;

	lut_sub lut_1816 ({sk[536], i_40_, i_39_, i_36_, i_37_, n_n515}, x1294x);
	defparam lut_1816.LUT_SIZE = 6;
	defparam lut_1816.mask = 64'h55ffffff00001040;

	lut_sub lut_1819 ({sk[537], i_39_, i_36_, i_38_}, n_n688);
	defparam lut_1819.LUT_SIZE = 4;
	defparam lut_1819.mask = 16'h1540;

	lut_sub lut_1821 ({sk[538], i_39_, i_36_, i_38_}, n_n918);
	defparam lut_1821.LUT_SIZE = 4;
	defparam lut_1821.mask = 16'h1508;

	lut_sub lut_1823 ({sk[539], i_16_, i_31_, x82x, n_n1066, x7288x, x7289x}, x726x);
	defparam lut_1823.LUT_SIZE = 7;
	defparam lut_1823.mask = 128'h77777f7f77777f7f07070000070f0000;

	lut_sub lut_1827 ({sk[540], i_16_, i_31_, n_n1066, x87x, x726x}, x725x);
	defparam lut_1827.LUT_SIZE = 6;
	defparam lut_1827.mask = 64'h55ffffff55555755;

	lut_sub lut_1830 ({sk[541], i_40_, i_39_, i_36_, i_35_, i_38_, x526x}, x1266x);
	defparam lut_1830.LUT_SIZE = 7;
	defparam lut_1830.mask = 128'h77777f7f77777f7f0000000000500010;

	lut_sub lut_1833 ({sk[542], i_7_, i_32_, i_34_, i_33_, i_35_}, x85x);
	defparam lut_1833.LUT_SIZE = 6;
	defparam lut_1833.mask = 64'h55ffffff20000000;

	lut_sub lut_1835 ({sk[543], i_40_, i_10_, i_27_, i_11_, i_36_, i_38_}, x7339x);
	defparam lut_1835.LUT_SIZE = 7;
	defparam lut_1835.mask = 128'h77777f7f77777f7f1111110020202020;

	lut_sub lut_1839 ({sk[544], i_40_, i_39_, i_38_, i_37_, n_n861, n_n991}, x1245x);
	defparam lut_1839.LUT_SIZE = 7;
	defparam lut_1839.mask = 128'h77777f7f77777f7f0001000111100000;

	lut_sub lut_1843 ({sk[545], i_34_, i_36_, i_35_, n_n861, n_n795, n_n977}, x7340x);
	defparam lut_1843.LUT_SIZE = 7;
	defparam lut_1843.mask = 128'h77777f7f77777f7f0003050000000000;

	lut_sub lut_1846 ({sk[546], i_40_, i_39_, i_36_, i_38_}, x371x);
	defparam lut_1846.LUT_SIZE = 5;
	defparam lut_1846.mask = 32'h00ff0080;

	lut_sub lut_1848 ({sk[547], i_24_, i_32_, x54x, x87x, n_n1023}, x245x);
	defparam lut_1848.LUT_SIZE = 6;
	defparam lut_1848.mask = 64'h55ffffff01000000;

	lut_sub lut_1850 ({sk[548], i_7_, i_5_, i_12_, i_11_, n_n848}, x364x);
	defparam lut_1850.LUT_SIZE = 6;
	defparam lut_1850.mask = 64'h55ffffff15000000;

	lut_sub lut_1853 ({sk[549], i_23_, i_32_, i_33_}, x7347x);
	defparam lut_1853.LUT_SIZE = 4;
	defparam lut_1853.mask = 16'h1540;

	lut_sub lut_1855 ({sk[550], i_40_, i_39_, i_35_, i_38_, n_n1074, x493x}, n_n857);
	defparam lut_1855.LUT_SIZE = 7;
	defparam lut_1855.mask = 128'h77777f7f77777f7f0000000000100000;

	lut_sub lut_1857 ({sk[551], i_9_, i_7_, i_5_}, n_n860);
	defparam lut_1857.LUT_SIZE = 4;
	defparam lut_1857.mask = 16'h1508;

	lut_sub lut_1859 ({sk[552], i_11_, i_18_, i_15_}, n_n859);
	defparam lut_1859.LUT_SIZE = 4;
	defparam lut_1859.mask = 16'h1501;

	lut_sub lut_1861 ({sk[553], i_12_, i_11_, i_18_, i_15_, i_19_}, x40x);
	defparam lut_1861.LUT_SIZE = 6;
	defparam lut_1861.mask = 64'h55ffffff00110313;

	lut_sub lut_1864 ({sk[554], i_9_, i_7_, i_5_, i_12_, i_11_, i_18_}, x44x);
	defparam lut_1864.LUT_SIZE = 7;
	defparam lut_1864.mask = 128'h77777f7f77777f7f150000001f000000;

	lut_sub lut_1868 ({sk[555], n_n1108, x155x, x7362x, x8561x}, n_n1577);
	defparam lut_1868.LUT_SIZE = 5;
	defparam lut_1868.mask = 32'h00ffbfff;

	lut_sub lut_1873 ({sk[556], i_2_, x314x, n_n926, n_n833, x7371x, x7367x}, n_n1575);
	defparam lut_1873.LUT_SIZE = 7;
	defparam lut_1873.mask = 128'h77777f7f77777f7f7777777777777fff;

	lut_sub lut_1878 ({sk[557], x181x, x431x, x79x, x149x, x318x, x1213x}, x7375x);
	defparam lut_1878.LUT_SIZE = 7;
	defparam lut_1878.mask = 128'h77777f7f77777f7f5f5f5f7fffffffff;

	lut_sub lut_1883 ({sk[558], n_n1118, n_n1113, x1675x, x6950x, x6951x, x7377x}, x7382x);
	defparam lut_1883.LUT_SIZE = 7;
	defparam lut_1883.mask = 128'h77777f7f77777f7f7fffffffffffffff;

	lut_sub lut_1890 ({sk[559], n_n979, x330x, n_n998, x60x, n_n791, x418x}, x641x);
	defparam lut_1890.LUT_SIZE = 7;
	defparam lut_1890.mask = 128'h77777f7f77777f7f0000557703035777;

	lut_sub lut_1894 ({sk[560], i_40_, n_n1001, x7347x, x360x, n_n843, x393x}, x7391x);
	defparam lut_1894.LUT_SIZE = 7;
	defparam lut_1894.mask = 128'h77777f7f77777f7f1111111f00000000;

	lut_sub lut_1897 ({sk[561], x406x, x60x, x321x, x360x, x7390x, x7389x}, x7392x);
	defparam lut_1897.LUT_SIZE = 7;
	defparam lut_1897.mask = 128'h77777f7f77777f7f0000030300550357;

	lut_sub lut_1900 ({sk[562], i_5_, i_11_, i_15_, i_34_, i_36_, i_35_}, x338x);
	defparam lut_1900.LUT_SIZE = 7;
	defparam lut_1900.mask = 128'h77777f7f77777f7f0000004000000000;

	lut_sub lut_1902 ({sk[563], i_40_, i_39_, i_38_, i_37_}, x60x);
	defparam lut_1902.LUT_SIZE = 5;
	defparam lut_1902.mask = 32'h00ff8040;

	lut_sub lut_1905 ({sk[564], i_22_, i_32_, i_33_}, x7406x);
	defparam lut_1905.LUT_SIZE = 4;
	defparam lut_1905.mask = 16'h1540;

	lut_sub lut_1907 ({sk[565], i_39_, n_n862, n_n488, x76x, x352x, x381x}, x1161x);
	defparam lut_1907.LUT_SIZE = 7;
	defparam lut_1907.mask = 128'h77777f7f77777f7f0000000000000057;

	lut_sub lut_1910 ({sk[566], i_21_, i_22_, x46x, x330x, n_n998, n_n949}, x1163x);
	defparam lut_1910.LUT_SIZE = 7;
	defparam lut_1910.mask = 128'h77777f7f77777f7f0001000100010000;

	lut_sub lut_1913 ({sk[567], i_40_, n_n1001, x7347x, x338x, x76x, x8573x}, x7429x);
	defparam lut_1913.LUT_SIZE = 7;
	defparam lut_1913.mask = 128'h77777f7f77777f7f2222222f22222222;

	lut_sub lut_1916 ({sk[568], i_3_, i_1_}, x675x);
	defparam lut_1916.LUT_SIZE = 3;
	defparam lut_1916.mask = 8'h37;

	lut_sub lut_1919 ({sk[569], i_3_, i_4_, i_1_, i_2_}, x677x);
	defparam lut_1919.LUT_SIZE = 5;
	defparam lut_1919.mask = 32'h00ff7fff;

	lut_sub lut_1924 ({sk[570], i_2_, n_n1055, n_n1001, x77x, x675x, x677x}, x7440x);
	defparam lut_1924.LUT_SIZE = 7;
	defparam lut_1924.mask = 128'h77777f7f77777f7f0005030700050f0f;

	lut_sub lut_1928 ({sk[571], i_40_, i_39_, i_36_, i_38_, i_37_}, x394x);
	defparam lut_1928.LUT_SIZE = 6;
	defparam lut_1928.mask = 64'h55ffffff00000100;

	lut_sub lut_1930 ({sk[572], i_4_, i_0_, i_32_, i_34_, i_33_, i_35_}, x332x);
	defparam lut_1930.LUT_SIZE = 7;
	defparam lut_1930.mask = 128'h77777f7f77777f7f0000000000002000;

	lut_sub lut_1932 ({sk[573], i_40_, i_9_, i_5_, i_39_, n_n862, x521x}, x8547x);
	defparam lut_1932.LUT_SIZE = 7;
	defparam lut_1932.mask = 128'h77777f7f77777f7fa8ffffffaaffffff;

	lut_sub lut_1946 ({sk[574], n_n1014, n_n1061, x76x, x394x, x332x, x8547x}, x7444x);
	defparam lut_1946.LUT_SIZE = 7;
	defparam lut_1946.mask = 128'h77777f7f77777f7f03ab03ab03ab33bb;

	lut_sub lut_1950 ({sk[575], i_39_, i_32_, i_33_, i_38_, i_37_, n_n998}, x384x);
	defparam lut_1950.LUT_SIZE = 7;
	defparam lut_1950.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_1952 ({sk[576], i_7_, i_5_, i_11_, i_21_, i_15_}, x365x);
	defparam lut_1952.LUT_SIZE = 6;
	defparam lut_1952.mask = 64'h55ffffff04000000;

	lut_sub lut_1954 ({sk[577], i_24_, i_22_, i_32_, i_34_, i_33_}, x476x);
	defparam lut_1954.LUT_SIZE = 6;
	defparam lut_1954.mask = 64'h55ffffff00004000;

	lut_sub lut_1956 ({sk[578], i_7_, i_5_, i_11_, i_15_, x476x}, n_n819);
	defparam lut_1956.LUT_SIZE = 6;
	defparam lut_1956.mask = 64'h55ffffff01000000;

	lut_sub lut_1958 ({sk[579], i_40_, i_39_, i_23_, i_24_, i_38_, x51x}, x475x);
	defparam lut_1958.LUT_SIZE = 7;
	defparam lut_1958.mask = 128'h77777f7f77777f7f0000010000000000;

	lut_sub lut_1960 ({sk[580], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x824x);
	defparam lut_1960.LUT_SIZE = 7;
	defparam lut_1960.mask = 128'h77777f7f77777f7f0800000004000000;

	lut_sub lut_1963 ({sk[581], n_n969, x329x, n_n819, x99x, n_n977, x386x}, x8522x);
	defparam lut_1963.LUT_SIZE = 7;
	defparam lut_1963.mask = 128'h77777f7f77777f7fffaafca8ffaaf0a0;

	lut_sub lut_1970 ({sk[582], x476x, x87x, x475x, x824x, x8522x}, x7455x);
	defparam lut_1970.LUT_SIZE = 6;
	defparam lut_1970.mask = 64'h55ffffffaaafaabf;

	lut_sub lut_1974 ({sk[583], i_7_, i_5_, i_12_, i_11_, i_15_, x476x}, x132x);
	defparam lut_1974.LUT_SIZE = 7;
	defparam lut_1974.mask = 128'h77777f7f77777f7f0111000000000000;

	lut_sub lut_1977 ({sk[584], i_24_, i_32_, i_34_, i_33_, n_n968}, x99x);
	defparam lut_1977.LUT_SIZE = 6;
	defparam lut_1977.mask = 64'h55ffffff00001000;

	lut_sub lut_1979 ({sk[585], i_40_, i_39_, i_38_}, n_n977);
	defparam lut_1979.LUT_SIZE = 4;
	defparam lut_1979.mask = 16'h1510;

	lut_sub lut_1981 ({sk[586], i_40_, i_39_, i_36_, i_38_, i_37_}, x718x);
	defparam lut_1981.LUT_SIZE = 6;
	defparam lut_1981.mask = 64'h55ffffffb0f0b0d0;

	lut_sub lut_1987 ({sk[587], i_9_, i_7_, i_17_, i_16_, x251x, x339x}, x7477x);
	defparam lut_1987.LUT_SIZE = 7;
	defparam lut_1987.mask = 128'h77777f7f77777f7f7773333373333333;

	lut_sub lut_1992 ({sk[588], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x356x);
	defparam lut_1992.LUT_SIZE = 7;
	defparam lut_1992.mask = 128'h77777f7f77777f7f2000000000000000;

	lut_sub lut_1994 ({sk[589], i_9_, i_7_, i_11_, x496x, x498x}, x1073x);
	defparam lut_1994.LUT_SIZE = 6;
	defparam lut_1994.mask = 64'h55ffffff00007030;

	lut_sub lut_1997 ({sk[590], i_36_, n_n1001, n_n980, x453x, x404x, x55x}, x1088x);
	defparam lut_1997.LUT_SIZE = 7;
	defparam lut_1997.mask = 128'h77777f7f77777f7f0000000700000000;

	lut_sub lut_2000 ({sk[591], i_7_, i_14_, i_12_, i_11_, n_n775, x351x}, x1089x);
	defparam lut_2000.LUT_SIZE = 7;
	defparam lut_2000.mask = 128'h77777f7f77777f7f1111111000000000;

	lut_sub lut_2004 ({sk[592], i_7_, n_n969, x51x, x61x, x394x, x428x}, x7485x);
	defparam lut_2004.LUT_SIZE = 7;
	defparam lut_2004.mask = 128'h77777f7f77777f7f111111f111111111;

	lut_sub lut_2007 ({sk[593], i_9_, i_7_, n_n1074, n_n977, n_n1073, x498x}, x691x);
	defparam lut_2007.LUT_SIZE = 7;
	defparam lut_2007.mask = 128'h77777f7f77777f7f0000000055570000;

	lut_sub lut_2010 ({sk[594], i_9_, i_7_, i_37_, n_n1011, n_n1047, x692x}, x1082x);
	defparam lut_2010.LUT_SIZE = 7;
	defparam lut_2010.mask = 128'h77777f7f77777f7f0000000000010000;

	lut_sub lut_2012 ({sk[595], i_7_, i_11_, n_n785, x351x, x67x, x1081x}, x1074x);
	defparam lut_2012.LUT_SIZE = 7;
	defparam lut_2012.mask = 128'h77777f7f77777f7f005f005700000000;

	lut_sub lut_2016 ({sk[596], i_9_, n_n833, x79x, x85x, x1071x, x792x}, x791x);
	defparam lut_2016.LUT_SIZE = 7;
	defparam lut_2016.mask = 128'h77777f7f77777f7f05370537053705ff;

	lut_sub lut_2020 ({sk[597], i_40_, i_39_, i_36_, i_38_, x392x, x428x}, x1061x);
	defparam lut_2020.LUT_SIZE = 7;
	defparam lut_2020.mask = 128'h77777f7f77777f7f3333373300000000;

	lut_sub lut_2023 ({sk[598], i_40_, n_n795, n_n1001, n_n983, n_n668, n_n976}, x7497x);
	defparam lut_2023.LUT_SIZE = 7;
	defparam lut_2023.mask = 128'h77777f7f77777f7f0003000300001111;

	lut_sub lut_2026 ({sk[599], i_36_, i_38_, i_37_}, n_n693);
	defparam lut_2026.LUT_SIZE = 4;
	defparam lut_2026.mask = 16'h1508;

	lut_sub lut_2028 ({sk[600], i_40_, i_7_, i_39_, i_11_, x45x, n_n693}, x182x);
	defparam lut_2028.LUT_SIZE = 7;
	defparam lut_2028.mask = 128'h77777f7f77777f7f0000000000010000;

	lut_sub lut_2030 ({sk[601], i_7_, i_5_, i_32_, n_n833, x371x, n_n1023}, x301x);
	defparam lut_2030.LUT_SIZE = 7;
	defparam lut_2030.mask = 128'h77777f7f77777f7f0000150000000000;

	lut_sub lut_2033 ({sk[602], i_9_, i_17_, i_16_}, x55x);
	defparam lut_2033.LUT_SIZE = 4;
	defparam lut_2033.mask = 16'h15c8;

	lut_sub lut_2036 ({sk[603], i_24_, i_22_, i_32_}, n_n428);
	defparam lut_2036.LUT_SIZE = 4;
	defparam lut_2036.mask = 16'h1502;

	lut_sub lut_2038 ({sk[604], i_40_, i_39_, i_36_, i_38_, i_37_, n_n1023}, x7513x);
	defparam lut_2038.LUT_SIZE = 7;
	defparam lut_2038.mask = 128'h77777f7f77777f7f0000000010000400;

	lut_sub lut_2041 ({sk[605], x82x, x101x, x87x, n_n1023, n_n428, x7513x}, x1038x);
	defparam lut_2041.LUT_SIZE = 7;
	defparam lut_2041.mask = 128'h77777f7f77777f7f0011001311111313;

	lut_sub lut_2046 ({sk[606], i_40_, i_39_, i_38_, x35x, n_n848, x77x}, x532x);
	defparam lut_2046.LUT_SIZE = 7;
	defparam lut_2046.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_2048 ({sk[607], i_36_, i_37_}, x493x);
	defparam lut_2048.LUT_SIZE = 3;
	defparam lut_2048.mask = 8'h34;

	lut_sub lut_2050 ({sk[608], i_39_, i_34_, i_36_, i_35_, i_38_, i_37_}, n_n775);
	defparam lut_2050.LUT_SIZE = 7;
	defparam lut_2050.mask = 128'h77777f7f77777f7f4000000000000000;

	lut_sub lut_2052 ({sk[609], i_12_, i_11_, i_31_, x46x, n_n775, x407x}, n_n2687);
	defparam lut_2052.LUT_SIZE = 7;
	defparam lut_2052.mask = 128'h77777f7f77777f7f0000010000000000;

	lut_sub lut_2054 ({sk[610], i_30_, i_32_, i_31_, i_34_, i_33_, i_35_}, x361x);
	defparam lut_2054.LUT_SIZE = 7;
	defparam lut_2054.mask = 128'h77777f7f77777f7f2000000000000000;

	lut_sub lut_2056 ({sk[611], i_9_, i_5_, i_12_, i_11_, i_15_}, x98x);
	defparam lut_2056.LUT_SIZE = 6;
	defparam lut_2056.mask = 64'h55ffffff00001000;

	lut_sub lut_2058 ({sk[612], i_9_, i_5_, i_12_, i_11_, i_15_}, x522x);
	defparam lut_2058.LUT_SIZE = 6;
	defparam lut_2058.mask = 64'h55ffffff00000400;

	lut_sub lut_2060 ({sk[613], i_40_, i_39_, i_38_}, n_n1072);
	defparam lut_2060.LUT_SIZE = 4;
	defparam lut_2060.mask = 16'h1501;

	lut_sub lut_2062 ({sk[614], i_5_, i_11_, i_15_}, n_n949);
	defparam lut_2062.LUT_SIZE = 4;
	defparam lut_2062.mask = 16'h1510;

	lut_sub lut_2064 ({sk[615], i_24_, i_21_, i_22_, i_32_, i_34_, i_33_}, x480x);
	defparam lut_2064.LUT_SIZE = 7;
	defparam lut_2064.mask = 128'h77777f7f77777f7f0000000000000040;

	lut_sub lut_2066 ({sk[616], i_5_, i_11_, i_15_, x480x}, n_n937);
	defparam lut_2066.LUT_SIZE = 5;
	defparam lut_2066.mask = 32'h00ff0100;

	lut_sub lut_2068 ({sk[617], i_23_, i_24_, i_22_, i_32_}, x7124x);
	defparam lut_2068.LUT_SIZE = 5;
	defparam lut_2068.mask = 32'h00ff0002;

	lut_sub lut_2070 ({sk[618], i_12_, i_11_, i_31_, x46x, n_n775, x407x}, x7535x);
	defparam lut_2070.LUT_SIZE = 7;
	defparam lut_2070.mask = 128'h77777f7f77777f7f0000010001000000;

	lut_sub lut_2073 ({sk[619], i_28_, i_29_, x361x, x457x, x140x}, x7536x);
	defparam lut_2073.LUT_SIZE = 6;
	defparam lut_2073.mask = 64'h55ffffff57555555;

	lut_sub lut_2076 ({sk[620], x480x, x386x, n_n947, x80x, x7145x, x7147x}, x7537x);
	defparam lut_2076.LUT_SIZE = 7;
	defparam lut_2076.mask = 128'h77777f7f77777f7f01010101010101ff;

	lut_sub lut_2079 ({sk[621], i_40_, i_39_, i_38_, x391x, x146x, x89x}, x8519x);
	defparam lut_2079.LUT_SIZE = 7;
	defparam lut_2079.mask = 128'h77777f7f77777f7fccccccc0ccc088cc;

	lut_sub lut_2090 ({sk[622], i_40_, i_39_, i_38_}, x120x);
	defparam lut_2090.LUT_SIZE = 4;
	defparam lut_2090.mask = 16'h1581;

	lut_sub lut_2093 ({sk[623], i_39_, i_23_, i_21_, i_38_, i_37_}, x7134x);
	defparam lut_2093.LUT_SIZE = 6;
	defparam lut_2093.mask = 64'h55ffffff00000002;

	lut_sub lut_2095 ({sk[624], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x386x);
	defparam lut_2095.LUT_SIZE = 7;
	defparam lut_2095.mask = 128'h77777f7f77777f7f0000000004000000;

	lut_sub lut_2097 ({sk[625], i_9_, i_5_, i_12_, i_11_}, x42x);
	defparam lut_2097.LUT_SIZE = 5;
	defparam lut_2097.mask = 32'h00ff0070;

	lut_sub lut_2100 ({sk[626], i_24_, i_22_, i_15_, n_n1074, n_n968, x42x}, x417x);
	defparam lut_2100.LUT_SIZE = 7;
	defparam lut_2100.mask = 128'h77777f7f77777f7f0000000000000001;

	lut_sub lut_2102 ({sk[627], i_5_, i_12_, i_15_}, n_n947);
	defparam lut_2102.LUT_SIZE = 4;
	defparam lut_2102.mask = 16'h1510;

	lut_sub lut_2104 ({sk[628], i_36_, i_35_, i_37_}, n_n1012);
	defparam lut_2104.LUT_SIZE = 4;
	defparam lut_2104.mask = 16'h1540;

	lut_sub lut_2106 ({sk[629], i_7_, i_3_, i_39_, i_4_, n_n985, x80x}, x7555x);
	defparam lut_2106.LUT_SIZE = 7;
	defparam lut_2106.mask = 128'h77777f7f77777f7f0100110000000000;

	lut_sub lut_2109 ({sk[630], n_n2793, x68x, x174x, x300x, x504x, x7577x}, n_n1283);
	defparam lut_2109.LUT_SIZE = 7;
	defparam lut_2109.mask = 128'h77777f7f77777f7f5fff7fffffffffff;

	lut_sub lut_2115 ({sk[631], x950x, x952x, x7582x, x7583x}, n_n1285);
	defparam lut_2115.LUT_SIZE = 5;
	defparam lut_2115.mask = 32'h00ff7fff;

	lut_sub lut_2120 ({sk[632], x356x, x367x, x6858x, x942x, x943x, x944x}, x7591x);
	defparam lut_2120.LUT_SIZE = 7;
	defparam lut_2120.mask = 128'h77777f7f77777f7f7f7f7f7f7f7f7fff;

	lut_sub lut_2125 ({sk[633], x7596x, x7597x, x7611x, x8518x}, x7614x);
	defparam lut_2125.LUT_SIZE = 5;
	defparam lut_2125.mask = 32'h00ffbfff;

	lut_sub lut_2130 ({sk[634], i_7_, i_11_, i_32_, i_36_, x325x, x322x}, x131x);
	defparam lut_2130.LUT_SIZE = 7;
	defparam lut_2130.mask = 128'h77777f7f77777f7f0000010000000000;

	lut_sub lut_2132 ({sk[635], i_40_, i_36_, i_35_, i_38_}, x402x);
	defparam lut_2132.LUT_SIZE = 5;
	defparam lut_2132.mask = 32'h00ff0004;

	lut_sub lut_2134 ({sk[636], i_40_, i_39_, i_36_, i_38_, i_37_, x315x}, x506x);
	defparam lut_2134.LUT_SIZE = 7;
	defparam lut_2134.mask = 128'h77777f7f77777f7f0000000000004000;

	lut_sub lut_2136 ({sk[637], i_12_, i_11_, x323x, x387x, n_n860, x321x}, x882x);
	defparam lut_2136.LUT_SIZE = 7;
	defparam lut_2136.mask = 128'h77777f7f77777f7f0013001300130003;

	lut_sub lut_2140 ({sk[638], i_39_, i_34_, i_35_, i_38_, i_37_, x106x}, x883x);
	defparam lut_2140.LUT_SIZE = 7;
	defparam lut_2140.mask = 128'h77777f7f77777f7f0040000000000000;

	lut_sub lut_2142 ({sk[639], i_37_, x66x, n_n964, x408x, x76x, x356x}, x884x);
	defparam lut_2142.LUT_SIZE = 7;
	defparam lut_2142.mask = 128'h77777f7f77777f7f0101010301010101;

	lut_sub lut_2145 ({sk[640], i_9_, i_7_, i_5_, n_n411, n_n859, x40x}, x8517x);
	defparam lut_2145.LUT_SIZE = 7;
	defparam lut_2145.mask = 128'h77777f7f77777f7ffffffffff8ffffff;

	lut_sub lut_2159 ({sk[641], i_15_, x90x, x491x, n_n880, x44x, x8517x}, x878x);
	defparam lut_2159.LUT_SIZE = 7;
	defparam lut_2159.mask = 128'h77777f7f77777f7f00000a0a00000a0b;

	lut_sub lut_2162 ({sk[642], i_23_, i_24_, i_32_, n_n833, x364x, n_n1023}, x130x);
	defparam lut_2162.LUT_SIZE = 7;
	defparam lut_2162.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_2164 ({sk[643], i_40_, i_38_, i_37_, x52x, n_n860, x86x}, x877x);
	defparam lut_2164.LUT_SIZE = 7;
	defparam lut_2164.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_2166 ({sk[644], i_4_, i_1_, i_0_}, n_n710);
	defparam lut_2166.LUT_SIZE = 4;
	defparam lut_2166.mask = 16'h1540;

	lut_sub lut_2168 ({sk[645], n_n1008, x50x, x85x, n_n528, x408x, x7652x}, x7655x);
	defparam lut_2168.LUT_SIZE = 7;
	defparam lut_2168.mask = 128'h77777f7f77777f7f0000030300550357;

	lut_sub lut_2171 ({sk[646], i_13_, n_n1064, x47x, n_n969, n_n888, n_n700}, x870x);
	defparam lut_2171.LUT_SIZE = 7;
	defparam lut_2171.mask = 128'h77777f7f77777f7f0001000100000011;

	lut_sub lut_2174 ({sk[647], i_37_, n_n979, n_n880, n_n960, x97x, x227x}, x7653x);
	defparam lut_2174.LUT_SIZE = 7;
	defparam lut_2174.mask = 128'h77777f7f77777f7f5555575755555577;

	lut_sub lut_2178 ({sk[648], i_7_, i_32_, i_34_, i_33_, i_36_, i_35_}, x499x);
	defparam lut_2178.LUT_SIZE = 7;
	defparam lut_2178.mask = 128'h77777f7f77777f7f0400000000000000;

	lut_sub lut_2180 ({sk[649], i_37_, n_n1021, n_n861, x358x, n_n883, n_n888}, x177x);
	defparam lut_2180.LUT_SIZE = 7;
	defparam lut_2180.mask = 128'h77777f7f77777f7f00110f1f00110011;

	lut_sub lut_2183 ({sk[650], i_40_, i_39_, i_38_, i_37_, x358x, x328x}, x7657x);
	defparam lut_2183.LUT_SIZE = 7;
	defparam lut_2183.mask = 128'h77777f7f77777f7f3000300030053000;

	lut_sub lut_2186 ({sk[651], i_30_, i_28_, i_29_, x47x, x361x, x321x}, x756x);
	defparam lut_2186.LUT_SIZE = 7;
	defparam lut_2186.mask = 128'h77777f7f77777f7f0503000705030507;

	lut_sub lut_2191 ({sk[652], i_24_, i_32_, i_33_, n_n853, n_n848}, n_n559);
	defparam lut_2191.LUT_SIZE = 6;
	defparam lut_2191.mask = 64'h55ffffff00000100;

	lut_sub lut_2193 ({sk[653], i_40_, i_22_, i_15_, n_n979, n_n945, x44x}, x507x);
	defparam lut_2193.LUT_SIZE = 7;
	defparam lut_2193.mask = 128'h77777f7f77777f7f0000000000000001;

	lut_sub lut_2195 ({sk[654], i_5_, i_12_, i_15_, i_34_, i_36_, i_35_}, x360x);
	defparam lut_2195.LUT_SIZE = 7;
	defparam lut_2195.mask = 128'h77777f7f77777f7f0000004000000000;

	lut_sub lut_2197 ({sk[655], i_22_, i_32_, i_33_}, x7390x);
	defparam lut_2197.LUT_SIZE = 4;
	defparam lut_2197.mask = 16'h1540;

	lut_sub lut_2199 ({sk[656], i_5_, i_22_, i_32_, i_33_, n_n979, x86x}, n_n164);
	defparam lut_2199.LUT_SIZE = 7;
	defparam lut_2199.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_2201 ({sk[657], i_24_, i_22_, x46x, n_n1001, x338x, x360x}, x446x);
	defparam lut_2201.LUT_SIZE = 7;
	defparam lut_2201.mask = 128'h77777f7f77777f7f0007000700050000;

	lut_sub lut_2205 ({sk[658], n_n977, n_n866, n_n888, x633x, x418x, x7694x}, x443x);
	defparam lut_2205.LUT_SIZE = 7;
	defparam lut_2205.mask = 128'h77777f7f77777f7f0000030300050307;

	lut_sub lut_2208 ({sk[659], n_n969, x360x, x7390x, n_n164, x446x, x443x}, n_n1195);
	defparam lut_2208.LUT_SIZE = 7;
	defparam lut_2208.mask = 128'h77777f7f77777f7f777777777f7f7fff;

	lut_sub lut_2213 ({sk[660], n_n979, n_n969, n_n949, n_n947, n_n791, x8515x}, x287x);
	defparam lut_2213.LUT_SIZE = 7;
	defparam lut_2213.mask = 128'h77777f7f77777f7f0222022202220323;

	lut_sub lut_2217 ({sk[661], i_9_, i_17_, i_16_, n_n1014, n_n1009, x7725x}, x282x);
	defparam lut_2217.LUT_SIZE = 7;
	defparam lut_2217.mask = 128'h77777f7f77777f7f0000000000010101;

	lut_sub lut_2220 ({sk[662], i_16_, x45x, x445x, n_n488, x421x, x7727x}, x283x);
	defparam lut_2220.LUT_SIZE = 7;
	defparam lut_2220.mask = 128'h77777f7f77777f7f0003050700000505;

	lut_sub lut_2223 ({sk[663], i_39_, i_22_, i_38_, i_37_, x46x, x338x}, x289x);
	defparam lut_2223.LUT_SIZE = 7;
	defparam lut_2223.mask = 128'h77777f7f77777f7f0000000000100000;

	lut_sub lut_2225 ({sk[664], x45x, n_n969, x338x, n_n488, n_n791, x8570x}, x7720x);
	defparam lut_2225.LUT_SIZE = 7;
	defparam lut_2225.mask = 128'h77777f7f77777f7f000000330a0a0a3b;

	lut_sub lut_2228 ({sk[665], i_5_, i_15_, n_n1074, x81x, x353x, x6739x}, n_n1203);
	defparam lut_2228.LUT_SIZE = 7;
	defparam lut_2228.mask = 128'h77777f7f77777f7f3075303000550000;

	lut_sub lut_2231 ({sk[666], i_40_, i_14_, i_38_, n_n1074, n_n970, x6739x}, x7733x);
	defparam lut_2231.LUT_SIZE = 7;
	defparam lut_2231.mask = 128'h77777f7f77777f7f0505000007050300;

	lut_sub lut_2234 ({sk[667], i_40_, i_39_, i_38_, x90x, x89x}, x7735x);
	defparam lut_2234.LUT_SIZE = 6;
	defparam lut_2234.mask = 64'h55ffffff35350035;

	lut_sub lut_2239 ({sk[668], i_3_, i_4_, o_15_, x384x, x427x, x664x}, x7737x);
	defparam lut_2239.LUT_SIZE = 7;
	defparam lut_2239.mask = 128'h77777f7f77777f7f11ff1fff1fff1fff;

	lut_sub lut_2244 ({sk[669], i_5_, i_39_, i_12_, x389x, x353x, x96x}, x8514x);
	defparam lut_2244.LUT_SIZE = 7;
	defparam lut_2244.mask = 128'h77777f7f77777f7faaff80c0aaffa0f0;

	lut_sub lut_2251 ({sk[670], i_40_, i_5_, i_39_, i_36_, i_38_}, x406x);
	defparam lut_2251.LUT_SIZE = 6;
	defparam lut_2251.mask = 64'h55ffffff00004000;

	lut_sub lut_2253 ({sk[671], i_30_, i_36_, x45x, n_n973, x406x, x347x}, x249x);
	defparam lut_2253.LUT_SIZE = 7;
	defparam lut_2253.mask = 128'h77777f7f77777f7f0000000500330037;

	lut_sub lut_2256 ({sk[672], i_28_, i_29_}, x202x);
	defparam lut_2256.LUT_SIZE = 3;
	defparam lut_2256.mask = 8'h37;

	lut_sub lut_2259 ({sk[673], i_3_, i_1_, i_0_, i_32_, n_n1066}, x69x);
	defparam lut_2259.LUT_SIZE = 6;
	defparam lut_2259.mask = 64'h55ffffff00040404;

	lut_sub lut_2262 ({sk[674], i_7_, i_5_, i_24_, i_15_, n_n978, x51x}, x189x);
	defparam lut_2262.LUT_SIZE = 7;
	defparam lut_2262.mask = 128'h77777f7f77777f7f1011000000000000;

	lut_sub lut_2265 ({sk[675], i_32_, n_n979, n_n462, x7019x, n_n1066, x8556x}, x7789x);
	defparam lut_2265.LUT_SIZE = 7;
	defparam lut_2265.mask = 128'h77777f7f77777f7f0003aaab0000aaaa;

	lut_sub lut_2268 ({sk[676], n_n861, n_n998, n_n977, n_n710, n_n799, n_n715}, x7790x);
	defparam lut_2268.LUT_SIZE = 7;
	defparam lut_2268.mask = 128'h77777f7f77777f7f0000000000050307;

	lut_sub lut_2271 ({sk[677], i_7_, i_32_, i_36_, i_38_, i_37_, n_n1023}, x439x);
	defparam lut_2271.LUT_SIZE = 7;
	defparam lut_2271.mask = 128'h77777f7f77777f7f0040000000000000;

	lut_sub lut_2273 ({sk[678], i_40_, i_34_, i_36_, i_35_, n_n861, n_n795}, x168x);
	defparam lut_2273.LUT_SIZE = 7;
	defparam lut_2273.mask = 128'h77777f7f77777f7f0000100001100000;

	lut_sub lut_2277 ({sk[679], i_40_, i_39_, i_38_, i_37_, x358x, x510x}, x7798x);
	defparam lut_2277.LUT_SIZE = 7;
	defparam lut_2277.mask = 128'h77777f7f77777f7f0050003000500000;

	lut_sub lut_2280 ({sk[680], x88x, n_n991, x6939x, n_n997, x339x, x7796x}, x7799x);
	defparam lut_2280.LUT_SIZE = 7;
	defparam lut_2280.mask = 128'h77777f7f77777f7f1111111111ff1fff;

	lut_sub lut_2284 ({sk[681], i_31_, n_n1074, x47x, x91x, x37x, x605x}, x147x);
	defparam lut_2284.LUT_SIZE = 7;
	defparam lut_2284.mask = 128'h77777f7f77777f7f00000000000c005d;

	lut_sub lut_2287 ({sk[682], i_37_, n_n979, n_n1008, n_n861, n_n883, x7803x}, x7810x);
	defparam lut_2287.LUT_SIZE = 7;
	defparam lut_2287.mask = 128'h77777f7f77777f7f010101010101010f;

	lut_sub lut_2290 ({sk[683], i_39_, i_17_, x85x, x7652x, n_n793, x353x}, x7812x);
	defparam lut_2290.LUT_SIZE = 7;
	defparam lut_2290.mask = 128'h77777f7f77777f7f111f000f11110000;

	lut_sub lut_2293 ({sk[684], i_24_, i_21_, i_22_, i_15_, i_32_}, x7006x);
	defparam lut_2293.LUT_SIZE = 6;
	defparam lut_2293.mask = 64'h55ffffff00000200;

	lut_sub lut_2295 ({sk[685], i_11_, x92x, x7006x, n_n860, n_n1023, x412x}, x129x);
	defparam lut_2295.LUT_SIZE = 7;
	defparam lut_2295.mask = 128'h77777f7f77777f7f0000001100000013;

	lut_sub lut_2298 ({sk[686], i_21_, x52x, n_n860, n_n859, x412x, x492x}, x136x);
	defparam lut_2298.LUT_SIZE = 7;
	defparam lut_2298.mask = 128'h77777f7f77777f7f0000111f00001111;

	lut_sub lut_2301 ({sk[687], i_9_, i_7_, i_5_, x52x, x70x}, x137x);
	defparam lut_2301.LUT_SIZE = 6;
	defparam lut_2301.mask = 64'h55ffffff00001000;

	lut_sub lut_2303 ({sk[688], i_17_, i_32_, i_33_}, n_n642);
	defparam lut_2303.LUT_SIZE = 4;
	defparam lut_2303.mask = 16'h1504;

	lut_sub lut_2305 ({sk[689], i_7_, i_5_, i_12_, i_11_, i_16_}, x114x);
	defparam lut_2305.LUT_SIZE = 6;
	defparam lut_2305.mask = 64'h55ffffff14000000;

	lut_sub lut_2308 ({sk[690], i_17_, i_16_, i_32_, i_33_}, x38x);
	defparam lut_2308.LUT_SIZE = 5;
	defparam lut_2308.mask = 32'h00ff0444;

	lut_sub lut_2311 ({sk[691], i_14_, i_12_, i_16_, i_15_, i_32_, i_33_}, x126x);
	defparam lut_2311.LUT_SIZE = 7;
	defparam lut_2311.mask = 128'h77777f7f77777f7f0000000400000000;

	lut_sub lut_2313 ({sk[692], i_34_, i_35_, i_37_}, n_n888);
	defparam lut_2313.LUT_SIZE = 4;
	defparam lut_2313.mask = 16'h1520;

	lut_sub lut_2315 ({sk[693], i_7_, i_5_, i_13_, i_12_, i_11_}, x408x);
	defparam lut_2315.LUT_SIZE = 6;
	defparam lut_2315.mask = 64'h55ffffff08000000;

	lut_sub lut_2317 ({sk[694], i_7_, i_5_, i_13_, i_15_, i_32_, i_33_}, x97x);
	defparam lut_2317.LUT_SIZE = 7;
	defparam lut_2317.mask = 128'h77777f7f77777f7f4000000000000000;

	lut_sub lut_2319 ({sk[695], i_40_, i_13_, i_36_, i_38_, x47x, x387x}, x227x);
	defparam lut_2319.LUT_SIZE = 7;
	defparam lut_2319.mask = 128'h77777f7f77777f7f0000000000001000;

	lut_sub lut_2321 ({sk[696], i_10_, i_27_, i_36_, i_38_, i_37_}, x7652x);
	defparam lut_2321.LUT_SIZE = 6;
	defparam lut_2321.mask = 64'h55ffffff02020200;

	lut_sub lut_2324 ({sk[697], i_9_, i_7_, i_5_, i_11_, i_15_}, x368x);
	defparam lut_2324.LUT_SIZE = 6;
	defparam lut_2324.mask = 64'h55ffffff10000000;

	lut_sub lut_2326 ({sk[698], i_16_, i_32_, i_31_, i_33_}, x6850x);
	defparam lut_2326.LUT_SIZE = 5;
	defparam lut_2326.mask = 32'h00ff4000;

	lut_sub lut_2328 ({sk[699], i_9_, i_7_, i_5_, i_12_, i_15_}, x367x);
	defparam lut_2328.LUT_SIZE = 6;
	defparam lut_2328.mask = 64'h55ffffff10000000;

	lut_sub lut_2330 ({sk[700], i_39_, i_23_, i_38_, x90x, x365x, n_n2456}, x7577x);
	defparam lut_2330.LUT_SIZE = 7;
	defparam lut_2330.mask = 128'h77777f7f77777f7f5755555555555555;

	lut_sub lut_2333 ({sk[701], i_40_, i_39_, i_36_, i_38_}, x7145x);
	defparam lut_2333.LUT_SIZE = 5;
	defparam lut_2333.mask = 32'h00ff0008;

	lut_sub lut_2335 ({sk[702], i_40_, i_39_, i_36_, i_38_, x80x}, x395x);
	defparam lut_2335.LUT_SIZE = 6;
	defparam lut_2335.mask = 64'h55ffffff00000040;

	lut_sub lut_2337 ({sk[703], i_40_, i_39_, i_36_, i_38_, i_37_}, x595x);
	defparam lut_2337.LUT_SIZE = 6;
	defparam lut_2337.mask = 64'h55ffffffc0004000;

	lut_sub lut_2340 ({sk[704], i_40_, i_39_, i_23_, i_38_, i_37_}, x7558x);
	defparam lut_2340.LUT_SIZE = 6;
	defparam lut_2340.mask = 64'h55ffffff00200000;

	lut_sub lut_2342 ({sk[705], i_22_, x82x, x50x, x87x, x595x, x7558x}, x7560x);
	defparam lut_2342.LUT_SIZE = 7;
	defparam lut_2342.mask = 128'h77777f7f77777f7f0007005700050055;

	lut_sub lut_2346 ({sk[706], i_22_, x82x, x50x, n_n833, x395x, x87x}, x8559x);
	defparam lut_2346.LUT_SIZE = 7;
	defparam lut_2346.mask = 128'h77777f7f77777f7feeeaccc8ffffffff;

	lut_sub lut_2352 ({sk[707], i_7_, i_5_, i_12_, i_11_}, x315x);
	defparam lut_2352.LUT_SIZE = 5;
	defparam lut_2352.mask = 32'h00ff8000;

	lut_sub lut_2354 ({sk[708], i_13_, i_12_, i_11_, i_32_, x47x, n_n1023}, n_n525);
	defparam lut_2354.LUT_SIZE = 7;
	defparam lut_2354.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_2356 ({sk[709], i_7_, i_36_, i_38_, i_37_, x80x, x464x}, x148x);
	defparam lut_2356.LUT_SIZE = 7;
	defparam lut_2356.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_2358 ({sk[710], i_39_, i_31_, i_38_, n_n1074, n_n1012, x408x}, x236x);
	defparam lut_2358.LUT_SIZE = 7;
	defparam lut_2358.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_2360 ({sk[711], i_40_, i_39_, i_36_, i_38_, i_37_}, x357x);
	defparam lut_2360.LUT_SIZE = 6;
	defparam lut_2360.mask = 64'h55ffffff20000000;

	lut_sub lut_2362 ({sk[712], i_40_, i_39_, i_38_, i_37_}, x441x);
	defparam lut_2362.LUT_SIZE = 5;
	defparam lut_2362.mask = 32'h00ff0010;

	lut_sub lut_2364 ({sk[713], x335x, n_n1064, x396x, n_n862, x76x, x6834x}, x7565x);
	defparam lut_2364.LUT_SIZE = 7;
	defparam lut_2364.mask = 128'h77777f7f77777f7f0000010100ff01ff;

	lut_sub lut_2367 ({sk[714], i_23_, x432x, x329x, x422x, x408x, x357x}, x7566x);
	defparam lut_2367.LUT_SIZE = 7;
	defparam lut_2367.mask = 128'h77777f7f77777f7f010101ff01010101;

	lut_sub lut_2370 ({sk[715], i_38_, x358x, x396x, n_n710, x441x, x89x}, x7567x);
	defparam lut_2370.LUT_SIZE = 7;
	defparam lut_2370.mask = 128'h77777f7f77777f7f0055035700000303;

	lut_sub lut_2373 ({sk[716], i_13_, n_n1064, x50x, n_n1052, x315x, x236x}, x7568x);
	defparam lut_2373.LUT_SIZE = 7;
	defparam lut_2373.mask = 128'h77777f7f77777f7f5555555755555555;

	lut_sub lut_2376 ({sk[717], i_32_, i_31_, i_34_, i_33_, i_36_, i_35_}, x353x);
	defparam lut_2376.LUT_SIZE = 7;
	defparam lut_2376.mask = 128'h77777f7f77777f7f0000080000000000;

	lut_sub lut_2378 ({sk[718], i_40_, i_16_, x313x, x6920x, n_n793, x353x}, x7775x);
	defparam lut_2378.LUT_SIZE = 7;
	defparam lut_2378.mask = 128'h77777f7f77777f7f111f000f11110000;

	lut_sub lut_2381 ({sk[719], i_7_, i_5_, x46x, x366x, x53x, x43x}, x212x);
	defparam lut_2381.LUT_SIZE = 7;
	defparam lut_2381.mask = 128'h77777f7f77777f7f0007000500050005;

	lut_sub lut_2384 ({sk[720], i_36_, i_35_, n_n973, x79x, x347x, x209x}, x7773x);
	defparam lut_2384.LUT_SIZE = 7;
	defparam lut_2384.mask = 128'h77777f7f77777f7f5555555555575555;

	lut_sub lut_2387 ({sk[721], i_36_, x81x, x50x, n_n975, x408x, n_n287}, x663x);
	defparam lut_2387.LUT_SIZE = 7;
	defparam lut_2387.mask = 128'h77777f7f77777f7f0505053705050505;

	lut_sub lut_2390 ({sk[722], i_39_, i_36_, x81x, x408x, x80x, x199x}, x7784x);
	defparam lut_2390.LUT_SIZE = 7;
	defparam lut_2390.mask = 128'h77777f7f77777f7f5555555555575555;

	lut_sub lut_2393 ({sk[723], i_13_, x45x, x325x, n_n1047, x97x, x506x}, x7785x);
	defparam lut_2393.LUT_SIZE = 7;
	defparam lut_2393.mask = 128'h77777f7f77777f7f0003555700030003;

	lut_sub lut_2396 ({sk[724], i_32_, x54x, n_n775, x463x, x408x, n_n1023}, x7786x);
	defparam lut_2396.LUT_SIZE = 7;
	defparam lut_2396.mask = 128'h77777f7f77777f7f000f111f000f000f;

	lut_sub lut_2399 ({sk[725], i_7_, i_32_, i_33_, n_n710, n_n715}, x398x);
	defparam lut_2399.LUT_SIZE = 6;
	defparam lut_2399.mask = 64'h55ffffff01000000;

	lut_sub lut_2401 ({sk[726], i_32_, i_34_, i_33_, i_36_, i_35_}, x91x);
	defparam lut_2401.LUT_SIZE = 6;
	defparam lut_2401.mask = 64'h55ffffff08000000;

	lut_sub lut_2403 ({sk[727], i_12_, i_11_, i_18_, i_15_, x359x, n_n1023}, x8560x);
	defparam lut_2403.LUT_SIZE = 7;
	defparam lut_2403.mask = 128'h77777f7f77777f7ffffffffefffefffe;

	lut_sub lut_2417 ({sk[728], i_9_, i_21_, i_19_, x47x, n_n428, x8560x}, x1791x);
	defparam lut_2417.LUT_SIZE = 7;
	defparam lut_2417.mask = 128'h77777f7f77777f7f0002000000000000;

	lut_sub lut_2419 ({sk[729], i_40_, i_39_, i_38_, i_37_}, x342x);
	defparam lut_2419.LUT_SIZE = 5;
	defparam lut_2419.mask = 32'h00ff0040;

	lut_sub lut_2421 ({sk[730], i_18_, i_21_, i_22_, n_n979, x86x, x70x}, x8550x);
	defparam lut_2421.LUT_SIZE = 7;
	defparam lut_2421.mask = 128'h77777f7f77777f7ffffafffafff8fffa;

	lut_sub lut_2435 ({sk[731], i_24_, i_32_, i_33_, n_n860, x342x, x8550x}, x1792x);
	defparam lut_2435.LUT_SIZE = 7;
	defparam lut_2435.mask = 128'h77777f7f77777f7f0000000000020000;

	lut_sub lut_2437 ({sk[732], i_12_, i_11_, i_18_, i_24_, i_22_, i_19_}, x8553x);
	defparam lut_2437.LUT_SIZE = 7;
	defparam lut_2437.mask = 128'h77777f7f77777f7ffffffcfdfcfffcfd;

	lut_sub lut_2453 ({sk[733], i_9_, i_21_, i_15_, x47x, n_n857, x8553x}, x1789x);
	defparam lut_2453.LUT_SIZE = 7;
	defparam lut_2453.mask = 128'h77777f7f77777f7f0002000000000000;

	lut_sub lut_2455 ({sk[734], i_36_, i_35_, i_37_}, n_n1073);
	defparam lut_2455.LUT_SIZE = 4;
	defparam lut_2455.mask = 16'h1580;

	lut_sub lut_2457 ({sk[735], i_36_, i_35_, i_38_}, n_n993);
	defparam lut_2457.LUT_SIZE = 4;
	defparam lut_2457.mask = 16'h1580;

	lut_sub lut_2459 ({sk[736], i_16_, i_31_, i_34_, i_33_, i_35_, x87x}, n_n535);
	defparam lut_2459.LUT_SIZE = 7;
	defparam lut_2459.mask = 128'h77777f7f77777f7f0000000004000000;

	lut_sub lut_2461 ({sk[737], i_9_, i_5_, i_11_}, n_n492);
	defparam lut_2461.LUT_SIZE = 4;
	defparam lut_2461.mask = 16'h1540;

	lut_sub lut_2463 ({sk[738], i_36_, i_38_, i_37_}, n_n1065);
	defparam lut_2463.LUT_SIZE = 4;
	defparam lut_2463.mask = 16'h1501;

	lut_sub lut_2465 ({sk[739], i_9_, i_5_, i_12_}, n_n488);
	defparam lut_2465.LUT_SIZE = 4;
	defparam lut_2465.mask = 16'h1540;

	lut_sub lut_2467 ({sk[740], i_3_, i_0_, i_32_}, n_n453);
	defparam lut_2467.LUT_SIZE = 4;
	defparam lut_2467.mask = 16'h1502;

	lut_sub lut_2469 ({sk[741], i_5_, i_15_}, x378x);
	defparam lut_2469.LUT_SIZE = 3;
	defparam lut_2469.mask = 8'h38;

	lut_sub lut_2471 ({sk[742], i_5_, i_13_, i_15_}, n_n884);
	defparam lut_2471.LUT_SIZE = 4;
	defparam lut_2471.mask = 16'h1580;

	lut_sub lut_2473 ({sk[743], i_9_, i_5_, i_11_, i_16_, i_15_}, x517x);
	defparam lut_2473.LUT_SIZE = 6;
	defparam lut_2473.mask = 64'h55ffffff04000000;

	lut_sub lut_2475 ({sk[744], i_40_, i_36_, i_35_, i_38_}, x401x);
	defparam lut_2475.LUT_SIZE = 5;
	defparam lut_2475.mask = 32'h00ff0080;

	lut_sub lut_2477 ({sk[745], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x103x);
	defparam lut_2477.LUT_SIZE = 7;
	defparam lut_2477.mask = 128'h77777f7f77777f7f0000a000c000e000;

	lut_sub lut_2480 ({sk[746], i_40_, i_5_, i_39_, i_36_, i_38_, i_37_}, x457x);
	defparam lut_2480.LUT_SIZE = 7;
	defparam lut_2480.mask = 128'h77777f7f77777f7f0040000000000000;

	lut_sub lut_2482 ({sk[747], i_5_, i_12_, i_17_, i_16_, i_15_}, x513x);
	defparam lut_2482.LUT_SIZE = 6;
	defparam lut_2482.mask = 64'h55ffffff00400000;

	lut_sub lut_2484 ({sk[748], i_21_, i_32_, i_33_}, n_n791);
	defparam lut_2484.LUT_SIZE = 4;
	defparam lut_2484.mask = 16'h1540;

	lut_sub lut_2486 ({sk[749], i_39_, n_n862, n_n492, x76x, x352x, x381x}, x1179x);
	defparam lut_2486.LUT_SIZE = 7;
	defparam lut_2486.mask = 128'h77777f7f77777f7f0000000000000057;

	lut_sub lut_2489 ({sk[750], i_30_, i_28_, i_29_, x361x, x457x, x321x}, x1181x);
	defparam lut_2489.LUT_SIZE = 7;
	defparam lut_2489.mask = 128'h77777f7f77777f7f0000030000110300;

	lut_sub lut_2492 ({sk[751], n_n560, x338x, x76x, x60x, x513x, n_n791}, x7417x);
	defparam lut_2492.LUT_SIZE = 7;
	defparam lut_2492.mask = 128'h77777f7f77777f7f0000050500330537;

	lut_sub lut_2495 ({sk[752], i_5_, i_31_, i_36_, i_35_}, x6739x);
	defparam lut_2495.LUT_SIZE = 5;
	defparam lut_2495.mask = 32'h00ff0800;

	lut_sub lut_2497 ({sk[753], i_5_, i_32_, i_31_, i_34_, i_33_, n_n964}, x96x);
	defparam lut_2497.LUT_SIZE = 7;
	defparam lut_2497.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_2499 ({sk[754], i_17_, i_16_, i_32_, i_31_, i_33_}, x6852x);
	defparam lut_2499.LUT_SIZE = 6;
	defparam lut_2499.mask = 64'h55ffffff40000000;

	lut_sub lut_2501 ({sk[755], i_40_, i_34_, i_36_, i_35_, i_38_, i_37_}, x1787x);
	defparam lut_2501.LUT_SIZE = 7;
	defparam lut_2501.mask = 128'h77777f7f77777f7f2000000000000000;

	lut_sub lut_2503 ({sk[756], i_40_, i_39_, i_34_, i_38_, i_37_, n_n964}, x64x);
	defparam lut_2503.LUT_SIZE = 7;
	defparam lut_2503.mask = 128'h77777f7f77777f7f1400040010000000;

	lut_sub lut_2506 ({sk[757], i_24_, i_32_, i_33_, n_n853, n_n850, n_n848}, x106x);
	defparam lut_2506.LUT_SIZE = 7;
	defparam lut_2506.mask = 128'h77777f7f77777f7f0000000000150000;

	lut_sub lut_2509 ({sk[758], i_32_, i_31_, i_34_, i_33_, i_35_}, x321x);
	defparam lut_2509.LUT_SIZE = 6;
	defparam lut_2509.mask = 64'h55ffffff20000000;

	lut_sub lut_2511 ({sk[759], i_21_, i_15_, i_19_, x90x, n_n978, x8552x}, x1780x);
	defparam lut_2511.LUT_SIZE = 7;
	defparam lut_2511.mask = 128'h77777f7f77777f7f0000020000000000;

	lut_sub lut_2513 ({sk[760], i_12_, i_17_, i_16_, x82x, n_n833, x321x}, x1781x);
	defparam lut_2513.LUT_SIZE = 7;
	defparam lut_2513.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_2515 ({sk[761], n_n1055, x94x, x368x, x6850x, x64x, x106x}, x8543x);
	defparam lut_2515.LUT_SIZE = 7;
	defparam lut_2515.mask = 128'h77777f7f77777f7ffffcfffcfffcaaa8;

	lut_sub lut_2525 ({sk[762], i_3_, i_4_, i_32_}, n_n1057);
	defparam lut_2525.LUT_SIZE = 4;
	defparam lut_2525.mask = 16'h1520;

	lut_sub lut_2527 ({sk[763], i_5_, i_24_, i_32_, i_33_, n_n979, x78x}, n_n459);
	defparam lut_2527.LUT_SIZE = 7;
	defparam lut_2527.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_2529 ({sk[764], i_5_, i_12_, i_11_}, n_n907);
	defparam lut_2529.LUT_SIZE = 4;
	defparam lut_2529.mask = 16'h1580;

	lut_sub lut_2531 ({sk[765], i_13_, i_34_, i_36_, i_35_, x46x, n_n907}, n_n905);
	defparam lut_2531.LUT_SIZE = 7;
	defparam lut_2531.mask = 128'h77777f7f77777f7f0100000000000000;

	lut_sub lut_2533 ({sk[766], i_38_, n_n1064, n_n1001, n_n836, n_n459, x524x}, x7402x);
	defparam lut_2533.LUT_SIZE = 7;
	defparam lut_2533.mask = 128'h77777f7f77777f7f0537373705370537;

	lut_sub lut_2537 ({sk[767], n_n1014, n_n1061, x69x, x154x, x394x, x426x}, x8525x);
	defparam lut_2537.LUT_SIZE = 7;
	defparam lut_2537.mask = 128'h77777f7f77777f7fe0e0e0e0e0e0a000;

	lut_sub lut_2543 ({sk[768], i_34_, i_36_, i_35_, i_37_}, x624x);
	defparam lut_2543.LUT_SIZE = 5;
	defparam lut_2543.mask = 32'h00ff1500;

	lut_sub lut_2546 ({sk[769], i_16_, i_15_}, x352x);
	defparam lut_2546.LUT_SIZE = 3;
	defparam lut_2546.mask = 8'h34;

	lut_sub lut_2548 ({sk[770], i_34_, i_33_, i_35_, n_n1057, n_n843}, x524x);
	defparam lut_2548.LUT_SIZE = 6;
	defparam lut_2548.mask = 64'h55ffffff00000010;

	lut_sub lut_2550 ({sk[771], i_9_, i_39_, i_11_, i_36_, i_38_, n_n947}, x8569x);
	defparam lut_2550.LUT_SIZE = 7;
	defparam lut_2550.mask = 128'h77777f7f77777f7fffffefffffffffff;

	lut_sub lut_2566 ({sk[772], i_16_, i_15_, i_36_, x81x, n_n488, x8569x}, x7713x);
	defparam lut_2566.LUT_SIZE = 7;
	defparam lut_2566.mask = 128'h77777f7f77777f7faaaaabaaaaaaaaaa;

	lut_sub lut_2569 ({sk[773], n_n880, x91x, n_n492, n_n488, x352x, x295x}, x7714x);
	defparam lut_2569.LUT_SIZE = 7;
	defparam lut_2569.mask = 128'h77777f7f77777f7f5555555555555777;

	lut_sub lut_2573 ({sk[774], i_40_, n_n836, n_n843, x518x, x524x, x383x}, x7715x);
	defparam lut_2573.LUT_SIZE = 7;
	defparam lut_2573.mask = 128'h77777f7f77777f7f111f333f000f333f;

	lut_sub lut_2577 ({sk[775], i_5_, i_12_, i_11_, i_15_, i_32_, i_33_}, x460x);
	defparam lut_2577.LUT_SIZE = 7;
	defparam lut_2577.mask = 128'h77777f7f77777f7f0004040000000000;

	lut_sub lut_2580 ({sk[776], i_22_, i_38_, i_37_, x46x, x338x, x360x}, x456x);
	defparam lut_2580.LUT_SIZE = 7;
	defparam lut_2580.mask = 128'h77777f7f77777f7f0007000000000000;

	lut_sub lut_2583 ({sk[777], i_24_, i_32_, i_33_, n_n1011, x338x, x360x}, x459x);
	defparam lut_2583.LUT_SIZE = 7;
	defparam lut_2583.mask = 128'h77777f7f77777f7f0007000000000000;

	lut_sub lut_2586 ({sk[778], x81x, n_n979, x323x, n_n791, x36x, x7687x}, x7691x);
	defparam lut_2586.LUT_SIZE = 7;
	defparam lut_2586.mask = 128'h77777f7f77777f7f0055005500550357;

	lut_sub lut_2589 ({sk[779], n_n960, n_n1073, x460x, x456x, x459x, x7691x}, n_n1193);
	defparam lut_2589.LUT_SIZE = 7;
	defparam lut_2589.mask = 128'h77777f7f77777f7f7f7f7f7f7f7f7fff;

	lut_sub lut_2594 ({sk[780], i_5_, i_12_, i_11_, i_15_}, x633x);
	defparam lut_2594.LUT_SIZE = 5;
	defparam lut_2594.mask = 32'h00ff1500;

	lut_sub lut_2597 ({sk[781], i_40_, i_10_, i_27_, i_39_, x45x, n_n1061}, x154x);
	defparam lut_2597.LUT_SIZE = 7;
	defparam lut_2597.mask = 128'h77777f7f77777f7f0000001000000000;

	lut_sub lut_2599 ({sk[782], i_40_, i_39_, i_32_, i_34_, i_33_}, x427x);
	defparam lut_2599.LUT_SIZE = 6;
	defparam lut_2599.mask = 64'h55ffffff00400000;

	lut_sub lut_2601 ({sk[783], i_9_, i_5_, i_12_, i_15_}, x635x);
	defparam lut_2601.LUT_SIZE = 5;
	defparam lut_2601.mask = 32'h00ffb000;

	lut_sub lut_2604 ({sk[784], i_40_, i_39_, i_36_, i_38_, i_37_, n_n874}, x233x);
	defparam lut_2604.LUT_SIZE = 7;
	defparam lut_2604.mask = 128'h77777f7f77777f7f0000000000001000;

	lut_sub lut_2606 ({sk[785], i_9_, i_7_, i_5_, i_12_, i_15_}, x7288x);
	defparam lut_2606.LUT_SIZE = 6;
	defparam lut_2606.mask = 64'h55ffffff00001000;

	lut_sub lut_2608 ({sk[786], i_16_, i_32_, i_31_, i_33_}, x6858x);
	defparam lut_2608.LUT_SIZE = 5;
	defparam lut_2608.mask = 32'h00ff4000;

	lut_sub lut_2610 ({sk[787], i_39_, i_17_, i_38_}, x6859x);
	defparam lut_2610.LUT_SIZE = 4;
	defparam lut_2610.mask = 16'h1504;

	lut_sub lut_2612 ({sk[788], i_34_, i_33_, i_36_, i_35_, n_n709, n_n1057}, x393x);
	defparam lut_2612.LUT_SIZE = 7;
	defparam lut_2612.mask = 128'h77777f7f77777f7f0000000000001000;

	lut_sub lut_2614 ({sk[789], i_30_, i_28_, i_29_}, x7389x);
	defparam lut_2614.LUT_SIZE = 4;
	defparam lut_2614.mask = 16'h1504;

	lut_sub lut_2616 ({sk[790], i_22_, i_32_, i_34_, i_33_, i_36_, i_35_}, x418x);
	defparam lut_2616.LUT_SIZE = 7;
	defparam lut_2616.mask = 128'h77777f7f77777f7f0008000000000000;

	lut_sub lut_2618 ({sk[791], i_9_, i_7_, i_5_, i_11_, i_17_, i_15_}, x6856x);
	defparam lut_2618.LUT_SIZE = 7;
	defparam lut_2618.mask = 128'h77777f7f77777f7f0400000000000000;

	lut_sub lut_2620 ({sk[792], i_39_, i_19_, i_38_, i_37_}, x6976x);
	defparam lut_2620.LUT_SIZE = 5;
	defparam lut_2620.mask = 32'h00ff4000;

	lut_sub lut_2622 ({sk[793], i_21_, i_32_, i_34_, i_33_, i_36_, i_35_}, x6977x);
	defparam lut_2622.LUT_SIZE = 7;
	defparam lut_2622.mask = 128'h77777f7f77777f7f0400000000000000;

	lut_sub lut_2624 ({sk[794], i_18_, i_21_, i_32_, i_33_, x368x}, n_n790);
	defparam lut_2624.LUT_SIZE = 6;
	defparam lut_2624.mask = 64'h55ffffff10000000;

	lut_sub lut_2626 ({sk[795], i_18_, n_n1055, n_n979, x368x, n_n791, x367x}, x950x);
	defparam lut_2626.LUT_SIZE = 7;
	defparam lut_2626.mask = 128'h77777f7f77777f7f0000001300000000;

	lut_sub lut_2629 ({sk[796], i_16_, i_31_, x46x, n_n775, x368x, x367x}, x952x);
	defparam lut_2629.LUT_SIZE = 7;
	defparam lut_2629.mask = 128'h77777f7f77777f7f0007000000000000;

	lut_sub lut_2632 ({sk[797], i_17_, i_31_, x46x, n_n775, x368x, x367x}, x7582x);
	defparam lut_2632.LUT_SIZE = 7;
	defparam lut_2632.mask = 128'h77777f7f77777f7f0007000000000000;

	lut_sub lut_2635 ({sk[798], x368x, x6850x, x356x, x367x, x6976x, x6977x}, x7583x);
	defparam lut_2635.LUT_SIZE = 7;
	defparam lut_2635.mask = 128'h77777f7f77777f7f01010101111111ff;

	lut_sub lut_2639 ({sk[799], i_7_, i_5_, i_12_, i_11_, i_15_}, x486x);
	defparam lut_2639.LUT_SIZE = 6;
	defparam lut_2639.mask = 64'h55ffffff15000000;

	lut_sub lut_2642 ({sk[800], i_17_, i_16_, i_32_, i_31_, i_33_, x82x}, n_n773);
	defparam lut_2642.LUT_SIZE = 7;
	defparam lut_2642.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_2644 ({sk[801], i_34_, i_36_, i_35_, i_37_, n_n880, n_n977}, x8515x);
	defparam lut_2644.LUT_SIZE = 7;
	defparam lut_2644.mask = 128'h77777f7f77777f7fffafffaffcffffff;

	lut_sub lut_2662 ({sk[802], i_17_, i_16_}, x110x);
	defparam lut_2662.LUT_SIZE = 3;
	defparam lut_2662.mask = 8'h3e;

	lut_sub lut_2665 ({sk[803], i_39_, i_32_, i_34_, i_33_, i_38_, n_n968}, x303x);
	defparam lut_2665.LUT_SIZE = 7;
	defparam lut_2665.mask = 128'h77777f7f77777f7f0000000001000000;

	lut_sub lut_2667 ({sk[804], i_40_, i_39_, i_32_, i_38_, i_37_, n_n976}, x331x);
	defparam lut_2667.LUT_SIZE = 7;
	defparam lut_2667.mask = 128'h77777f7f77777f7f0400000000000000;

	lut_sub lut_2669 ({sk[805], i_14_, i_12_, i_11_, i_32_, i_33_, i_35_}, x7725x);
	defparam lut_2669.LUT_SIZE = 7;
	defparam lut_2669.mask = 128'h77777f7f77777f7f0000000000000020;

	lut_sub lut_2671 ({sk[806], i_39_, i_17_, i_36_, i_38_, i_37_}, x7727x);
	defparam lut_2671.LUT_SIZE = 6;
	defparam lut_2671.mask = 64'h55ffffff40000000;

	lut_sub lut_2673 ({sk[807], i_40_, i_39_, i_32_, i_34_, i_33_}, x6826x);
	defparam lut_2673.LUT_SIZE = 6;
	defparam lut_2673.mask = 64'h55ffffff00000010;

	lut_sub lut_2675 ({sk[808], i_40_, i_39_, i_36_, i_35_, i_38_, n_n966}, x336x);
	defparam lut_2675.LUT_SIZE = 7;
	defparam lut_2675.mask = 128'h77777f7f77777f7f0000000000004000;

	lut_sub lut_2677 ({sk[809], i_2_, i_0_, i_32_}, n_n458);
	defparam lut_2677.LUT_SIZE = 4;
	defparam lut_2677.mask = 16'h1502;

	lut_sub lut_2679 ({sk[810], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x7468x);
	defparam lut_2679.LUT_SIZE = 7;
	defparam lut_2679.mask = 128'h77777f7f77777f7f00008000c400a200;

	lut_sub lut_2684 ({sk[811], i_2_, i_0_, i_32_, i_34_, i_33_, i_35_}, x426x);
	defparam lut_2684.LUT_SIZE = 7;
	defparam lut_2684.mask = 128'h77777f7f77777f7f0000000000002000;

	lut_sub lut_2686 ({sk[812], i_17_, i_16_, i_32_, i_33_}, x351x);
	defparam lut_2686.LUT_SIZE = 5;
	defparam lut_2686.mask = 32'h00ff0004;

	lut_sub lut_2688 ({sk[813], i_40_, i_38_}, x343x);
	defparam lut_2688.LUT_SIZE = 3;
	defparam lut_2688.mask = 8'h34;

	lut_sub lut_2690 ({sk[814], i_5_, i_35_, i_38_, i_37_}, x664x);
	defparam lut_2690.LUT_SIZE = 5;
	defparam lut_2690.mask = 32'h00ff4404;

	lut_sub lut_2693 ({sk[815], i_32_, i_34_, i_33_, i_36_, i_35_}, x397x);
	defparam lut_2693.LUT_SIZE = 6;
	defparam lut_2693.mask = 64'h55ffffff02000000;

	lut_sub lut_2695 ({sk[816], i_10_, i_39_, i_38_, i_37_, x46x, n_n991}, x184x);
	defparam lut_2695.LUT_SIZE = 7;
	defparam lut_2695.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_2697 ({sk[817], i_27_, i_39_, i_38_, i_37_, x46x, n_n991}, x187x);
	defparam lut_2697.LUT_SIZE = 7;
	defparam lut_2697.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_2699 ({sk[818], i_30_, i_29_}, x53x);
	defparam lut_2699.LUT_SIZE = 3;
	defparam lut_2699.mask = 8'h36;

	lut_sub lut_2702 ({sk[819], i_12_, i_11_}, x41x);
	defparam lut_2702.LUT_SIZE = 3;
	defparam lut_2702.mask = 8'h3e;

	lut_sub lut_2705 ({sk[820], x50x, x54x, x371x, x408x, x76x, x103x}, x6861x);
	defparam lut_2705.LUT_SIZE = 7;
	defparam lut_2705.mask = 128'h77777f7f77777f7f01010101010f0f0f;

	lut_sub lut_2709 ({sk[821], i_14_, i_12_}, x67x);
	defparam lut_2709.LUT_SIZE = 3;
	defparam lut_2709.mask = 8'h3e;

	lut_sub lut_2712 ({sk[822], i_40_, i_38_, i_37_}, x403x);
	defparam lut_2712.LUT_SIZE = 4;
	defparam lut_2712.mask = 16'h1540;

	lut_sub lut_2714 ({sk[823], i_3_, i_1_, i_2_, i_0_, i_32_, n_n1023}, x680x);
	defparam lut_2714.LUT_SIZE = 7;
	defparam lut_2714.mask = 128'h77777f7f77777f7f0404000404040404;

	lut_sub lut_2718 ({sk[824], i_39_, i_36_, i_35_, i_38_, i_37_}, x521x);
	defparam lut_2718.LUT_SIZE = 6;
	defparam lut_2718.mask = 64'h55ffffff00001000;

	lut_sub lut_2720 ({sk[825], i_0_, i_32_, i_33_, i_37_, n_n979}, x413x);
	defparam lut_2720.LUT_SIZE = 6;
	defparam lut_2720.mask = 64'h55ffffff00000100;

	lut_sub lut_2722 ({sk[826], i_1_, i_0_}, x318x);
	defparam lut_2722.LUT_SIZE = 3;
	defparam lut_2722.mask = 8'h31;

	lut_sub lut_2724 ({sk[827], i_32_, n_n1066, n_n453, n_n458, x332x, x318x}, x683x);
	defparam lut_2724.LUT_SIZE = 7;
	defparam lut_2724.mask = 128'h77777f7f77777f7f33337fff33333fff;

	lut_sub lut_2729 ({sk[828], i_12_, i_11_, i_18_, i_15_, n_n793, x303x}, x1765x);
	defparam lut_2729.LUT_SIZE = 7;
	defparam lut_2729.mask = 128'h77777f7f77777f7f0000010001000100;

	lut_sub lut_2732 ({sk[829], i_40_, i_38_, i_37_, n_n964, x408x, x76x}, x1766x);
	defparam lut_2732.LUT_SIZE = 7;
	defparam lut_2732.mask = 128'h77777f7f77777f7f0000010000000000;

	lut_sub lut_2734 ({sk[830], i_31_, n_n1074, n_n1012, n_n2456, n_n799, x6862x}, x6868x);
	defparam lut_2734.LUT_SIZE = 7;
	defparam lut_2734.mask = 128'h77777f7f77777f7f0f0f0f1f0f0f0f0f;

	lut_sub lut_2737 ({sk[831], i_40_, i_39_, i_36_, i_38_, i_37_}, x710x);
	defparam lut_2737.LUT_SIZE = 6;
	defparam lut_2737.mask = 64'h55ffffff8020c020;

	lut_sub lut_2741 ({sk[832], i_24_, i_32_, x82x, n_n1023, x710x}, n_n1113);
	defparam lut_2741.LUT_SIZE = 6;
	defparam lut_2741.mask = 64'h55ffffff01000000;

	lut_sub lut_2743 ({sk[833], i_21_, x82x, x50x, n_n833, x87x, n_n1113}, x6877x);
	defparam lut_2743.LUT_SIZE = 7;
	defparam lut_2743.mask = 128'h77777f7f77777f7f555555555557555f;

	lut_sub lut_2747 ({sk[834], n_n979, n_n158, n_n853, n_n850, n_n469, x304x}, x1751x);
	defparam lut_2747.LUT_SIZE = 7;
	defparam lut_2747.mask = 128'h77777f7f77777f7f0000000000000777;

	lut_sub lut_2752 ({sk[835], x93x, n_n469, x371x, n_n834, n_n527, x246x}, x8562x);
	defparam lut_2752.LUT_SIZE = 7;
	defparam lut_2752.mask = 128'h77777f7f77777f7ffff0aaa0fff08880;

	lut_sub lut_2759 ({sk[836], i_7_, i_3_, i_4_, i_0_, n_n1074, x431x}, x149x);
	defparam lut_2759.LUT_SIZE = 7;
	defparam lut_2759.mask = 128'h77777f7f77777f7f0001010100000000;

	lut_sub lut_2762 ({sk[837], i_7_, i_3_, i_4_, i_0_, n_n1074, x362x}, x155x);
	defparam lut_2762.LUT_SIZE = 7;
	defparam lut_2762.mask = 128'h77777f7f77777f7f0001010100000000;

	lut_sub lut_2765 ({sk[838], i_39_, n_n330, x385x, x387x, x65x, x383x}, x6892x);
	defparam lut_2765.LUT_SIZE = 7;
	defparam lut_2765.mask = 128'h77777f7f77777f7f0033003300330537;

	lut_sub lut_2768 ({sk[839], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x711x);
	defparam lut_2768.LUT_SIZE = 7;
	defparam lut_2768.mask = 128'h77777f7f77777f7f0000000000100020;

	lut_sub lut_2771 ({sk[840], i_38_, n_n1008, x429x, x79x, x711x, x6895x}, n_n1108);
	defparam lut_2771.LUT_SIZE = 7;
	defparam lut_2771.mask = 128'h77777f7f77777f7f0033003300330537;

	lut_sub lut_2774 ({sk[841], i_30_, i_7_, i_5_, i_28_, i_29_}, x689x);
	defparam lut_2774.LUT_SIZE = 6;
	defparam lut_2774.mask = 64'h55ffffff20004000;

	lut_sub lut_2777 ({sk[842], i_40_, i_7_, i_5_, i_15_, x93x, n_n1001}, x1731x);
	defparam lut_2777.LUT_SIZE = 7;
	defparam lut_2777.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_2779 ({sk[843], x313x, x422x, n_n462, n_n1065, x464x, x689x}, x6901x);
	defparam lut_2779.LUT_SIZE = 7;
	defparam lut_2779.mask = 128'h77777f7f77777f7f0000005503030357;

	lut_sub lut_2782 ({sk[844], i_16_, i_32_, i_31_}, n_n927);
	defparam lut_2782.LUT_SIZE = 4;
	defparam lut_2782.mask = 16'h1508;

	lut_sub lut_2784 ({sk[845], i_9_, i_7_}, x344x);
	defparam lut_2784.LUT_SIZE = 3;
	defparam lut_2784.mask = 8'h32;

	lut_sub lut_2786 ({sk[846], i_14_, i_12_, i_11_, i_17_, i_16_, x46x}, x692x);
	defparam lut_2786.LUT_SIZE = 7;
	defparam lut_2786.mask = 128'h77777f7f77777f7f1515151515151500;

	lut_sub lut_2793 ({sk[847], i_39_, i_34_, i_38_, i_37_, n_n964, x38x}, x498x);
	defparam lut_2793.LUT_SIZE = 7;
	defparam lut_2793.mask = 128'h77777f7f77777f7f0000000000100000;

	lut_sub lut_2795 ({sk[848], i_17_, i_16_, i_15_, n_n949, n_n492, x76x}, x7426x);
	defparam lut_2795.LUT_SIZE = 7;
	defparam lut_2795.mask = 128'h77777f7f77777f7f0515001100110000;

	lut_sub lut_2799 ({sk[849], i_7_, i_5_, i_28_, i_29_}, x43x);
	defparam lut_2799.LUT_SIZE = 5;
	defparam lut_2799.mask = 32'h00ff9000;

	lut_sub lut_2802 ({sk[850], i_30_, i_7_, i_5_, i_28_, i_29_}, x102x);
	defparam lut_2802.LUT_SIZE = 6;
	defparam lut_2802.mask = 64'h55ffffff9000b000;

	lut_sub lut_2806 ({sk[851], x330x, n_n998, n_n330, x387x, x97x, x119x}, x7663x);
	defparam lut_2806.LUT_SIZE = 7;
	defparam lut_2806.mask = 128'h77777f7f77777f7f0005000500053337;

	lut_sub lut_2809 ({sk[852], i_7_, i_5_, i_12_, i_34_, n_n964, n_n1048}, x246x);
	defparam lut_2809.LUT_SIZE = 7;
	defparam lut_2809.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_2811 ({sk[853], i_18_, i_21_, i_32_, i_33_}, x6968x);
	defparam lut_2811.LUT_SIZE = 5;
	defparam lut_2811.mask = 32'h00ff4000;

	lut_sub lut_2813 ({sk[854], i_7_, i_32_}, x376x);
	defparam lut_2813.LUT_SIZE = 3;
	defparam lut_2813.mask = 8'h38;

	lut_sub lut_2815 ({sk[855], i_7_, i_14_, i_15_, x322x, x110x, x41x}, n_n550);
	defparam lut_2815.LUT_SIZE = 7;
	defparam lut_2815.mask = 128'h77777f7f77777f7f0000000800000000;

	lut_sub lut_2817 ({sk[856], i_40_, i_39_, i_13_, x80x, x315x, x321x}, x854x);
	defparam lut_2817.LUT_SIZE = 7;
	defparam lut_2817.mask = 128'h77777f7f77777f7f0000000011110300;

	lut_sub lut_2820 ({sk[857], i_13_, i_12_, n_n527, x76x, x401x, x8572x}, x7667x);
	defparam lut_2820.LUT_SIZE = 7;
	defparam lut_2820.mask = 128'h77777f7f77777f7f00aa000000ab0000;

	lut_sub lut_2823 ({sk[858], n_n515, n_n330, x92x, x387x, x236x, x357x}, x8516x);
	defparam lut_2823.LUT_SIZE = 7;
	defparam lut_2823.mask = 128'h77777f7f77777f7fccccc8c8cc00c800;

	lut_sub lut_2830 ({sk[859], i_21_, i_15_, i_19_}, x492x);
	defparam lut_2830.LUT_SIZE = 4;
	defparam lut_2830.mask = 16'h1510;

	lut_sub lut_2832 ({sk[860], i_12_, i_11_, i_18_, i_21_, i_15_, i_19_}, x70x);
	defparam lut_2832.LUT_SIZE = 7;
	defparam lut_2832.mask = 128'h77777f7f77777f7f0000101010301030;

	lut_sub lut_2836 ({sk[861], i_36_, i_37_}, x383x);
	defparam lut_2836.LUT_SIZE = 3;
	defparam lut_2836.mask = 8'h38;

	lut_sub lut_2838 ({sk[862], i_38_, n_n842, x541x, x362x, x502x, n_n843}, x7362x);
	defparam lut_2838.LUT_SIZE = 7;
	defparam lut_2838.mask = 128'h77777f7f77777f7f000f000f000f111f;

	lut_sub lut_2841 ({sk[863], i_39_, x396x, n_n966, x371x, n_n834, n_n993}, x8561x);
	defparam lut_2841.LUT_SIZE = 7;
	defparam lut_2841.mask = 128'h77777f7f77777f7ffcfcfca8fcfcfcfc;

	lut_sub lut_2850 ({sk[864], i_7_, i_39_, i_32_, i_36_, i_38_, n_n1066}, x1109x);
	defparam lut_2850.LUT_SIZE = 7;
	defparam lut_2850.mask = 128'h77777f7f77777f7f4000000000000000;

	lut_sub lut_2852 ({sk[865], i_39_, i_34_, i_33_, i_36_, i_38_, i_37_}, x1110x);
	defparam lut_2852.LUT_SIZE = 7;
	defparam lut_2852.mask = 128'h77777f7f77777f7f0040000000200000;

	lut_sub lut_2855 ({sk[866], i_40_, i_34_, i_36_, i_35_, i_38_, i_37_}, x139x);
	defparam lut_2855.LUT_SIZE = 7;
	defparam lut_2855.mask = 128'h77777f7f77777f7f0400000007000000;

	lut_sub lut_2858 ({sk[867], i_9_, i_7_, i_15_, i_34_, i_33_, x8549x}, x1277x);
	defparam lut_2858.LUT_SIZE = 7;
	defparam lut_2858.mask = 128'h77777f7f77777f7f0000000000100000;

	lut_sub lut_2860 ({sk[868], i_31_, i_33_}, x488x);
	defparam lut_2860.LUT_SIZE = 3;
	defparam lut_2860.mask = 8'h34;

	lut_sub lut_2862 ({sk[869], i_39_, i_34_, i_35_, i_38_, i_37_}, x7317x);
	defparam lut_2862.LUT_SIZE = 6;
	defparam lut_2862.mask = 64'h55ffffff08000000;

	lut_sub lut_2864 ({sk[870], n_n853, n_n850, n_n945, n_n848, x139x, x7317x}, x7321x);
	defparam lut_2864.LUT_SIZE = 7;
	defparam lut_2864.mask = 128'h77777f7f77777f7f0000000700050007;

	lut_sub lut_2868 ({sk[871], i_38_, n_n964, n_n860, x166x, x1273x, x7314x}, x7319x);
	defparam lut_2868.LUT_SIZE = 7;
	defparam lut_2868.mask = 128'h77777f7f77777f7f3333333333333373;

	lut_sub lut_2871 ({sk[872], i_9_, i_7_, i_5_, i_11_, i_15_}, x7289x);
	defparam lut_2871.LUT_SIZE = 6;
	defparam lut_2871.mask = 64'h55ffffff00001000;

	lut_sub lut_2873 ({sk[873], i_12_, i_11_, i_16_, i_15_, i_32_, i_31_}, x1633x);
	defparam lut_2873.LUT_SIZE = 7;
	defparam lut_2873.mask = 128'h77777f7f77777f7f0000000800000000;

	lut_sub lut_2875 ({sk[874], i_40_, i_39_, i_32_, n_n985, n_n1009, n_n1023}, x1047x);
	defparam lut_2875.LUT_SIZE = 7;
	defparam lut_2875.mask = 128'h77777f7f77777f7f0000000005001100;

	lut_sub lut_2878 ({sk[875], i_2_, x314x, n_n833, x79x, x346x, x6895x}, x7605x);
	defparam lut_2878.LUT_SIZE = 7;
	defparam lut_2878.mask = 128'h77777f7f77777f7f01010101010101ff;

	lut_sub lut_2881 ({sk[876], i_9_, i_14_, i_17_, i_16_, i_32_, i_33_}, x1081x);
	defparam lut_2881.LUT_SIZE = 7;
	defparam lut_2881.mask = 128'h77777f7f77777f7f0000000004440000;

	lut_sub lut_2884 ({sk[877], i_40_, i_7_, i_39_, i_38_, n_n1074, n_n1073}, x496x);
	defparam lut_2884.LUT_SIZE = 7;
	defparam lut_2884.mask = 128'h77777f7f77777f7f0001000000000000;

	lut_sub lut_2886 ({sk[878], i_25_, n_n709, x324x, n_n969, n_n971, n_n966}, x6740x);
	defparam lut_2886.LUT_SIZE = 7;
	defparam lut_2886.mask = 128'h77777f7f77777f7f01010101010101ff;

	lut_sub lut_2889 ({sk[879], i_12_, i_15_, x90x, n_n967, x89x, x96x}, x6741x);
	defparam lut_2889.LUT_SIZE = 7;
	defparam lut_2889.mask = 128'h77777f7f77777f7f575f575f575f030f;

	lut_sub lut_2894 ({sk[880], i_40_, i_39_, i_38_, n_n1074, n_n968, n_n1073}, x6745x);
	defparam lut_2894.LUT_SIZE = 7;
	defparam lut_2894.mask = 128'h77777f7f77777f7f0300050007000505;

	lut_sub lut_2899 ({sk[881], i_40_, i_39_, i_38_, i_37_}, x124x);
	defparam lut_2899.LUT_SIZE = 5;
	defparam lut_2899.mask = 32'h00ff0888;

	lut_sub lut_2902 ({sk[882], i_12_, i_11_, i_15_}, x166x);
	defparam lut_2902.LUT_SIZE = 4;
	defparam lut_2902.mask = 16'h15fe;

	lut_sub lut_2906 ({sk[883], i_40_, i_39_, i_17_, i_16_, i_38_, i_37_}, x750x);
	defparam lut_2906.LUT_SIZE = 7;
	defparam lut_2906.mask = 128'h77777f7f77777f7ffbbbfffffbbbfddd;

	lut_sub lut_2913 ({sk[884], i_39_, i_34_, i_36_, i_35_, i_38_, i_37_}, x7334x);
	defparam lut_2913.LUT_SIZE = 7;
	defparam lut_2913.mask = 128'h77777f7f77777f7f0008000000580000;

	lut_sub lut_2916 ({sk[885], i_30_, i_32_, i_31_, x202x, n_n976, x458x}, x140x);
	defparam lut_2916.LUT_SIZE = 7;
	defparam lut_2916.mask = 128'h77777f7f77777f7f1000000000000000;

	lut_sub lut_2918 ({sk[886], i_5_, i_12_, i_11_, i_21_, i_22_, i_15_}, x7147x);
	defparam lut_2918.LUT_SIZE = 7;
	defparam lut_2918.mask = 128'h77777f7f77777f7f0001010100000000;

	lut_sub lut_2921 ({sk[887], i_7_, i_5_, i_29_}, x494x);
	defparam lut_2921.LUT_SIZE = 4;
	defparam lut_2921.mask = 16'h1540;

	lut_sub lut_2923 ({sk[888], i_21_, i_15_, i_32_, n_n853, n_n1023}, n_n765);
	defparam lut_2923.LUT_SIZE = 6;
	defparam lut_2923.mask = 64'h55ffffff00100000;

	lut_sub lut_2925 ({sk[889], i_30_, i_7_, i_5_, i_28_, i_29_}, x765x);
	defparam lut_2925.LUT_SIZE = 6;
	defparam lut_2925.mask = 64'h55ffffffd000b000;

	lut_sub lut_2930 ({sk[890], i_32_, i_34_, i_33_, i_36_, i_35_, i_37_}, x770x);
	defparam lut_2930.LUT_SIZE = 7;
	defparam lut_2930.mask = 128'h77777f7f77777f7f0021008000000000;

	lut_sub lut_2934 ({sk[891], i_40_, i_39_, i_38_, x389x, x51x, x770x}, x7162x);
	defparam lut_2934.LUT_SIZE = 7;
	defparam lut_2934.mask = 128'h77777f7f77777f7f0f33000000005500;

	lut_sub lut_2938 ({sk[892], i_3_, i_4_, i_1_, x314x, n_n926, n_n833}, x7371x);
	defparam lut_2938.LUT_SIZE = 7;
	defparam lut_2938.mask = 128'h77777f7f77777f7f0005050507070707;

	lut_sub lut_2943 ({sk[893], i_1_, o_32_, x88x, x314x, x6811x, n_n926}, x7367x);
	defparam lut_2943.LUT_SIZE = 7;
	defparam lut_2943.mask = 128'h77777f7f77777f7f0033ffff0537ffff;

	lut_sub lut_2947 ({sk[894], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x775x);
	defparam lut_2947.LUT_SIZE = 7;
	defparam lut_2947.mask = 128'h77777f7f77777f7f0808000000000a00;

	lut_sub lut_2950 ({sk[895], i_24_, i_22_, n_n1014, x51x, x417x, x380x}, x1489x);
	defparam lut_2950.LUT_SIZE = 7;
	defparam lut_2950.mask = 128'h77777f7f77777f7f0033003300330037;

	lut_sub lut_2953 ({sk[896], i_5_, x480x, x386x, x86x, x78x, x775x}, x7129x);
	defparam lut_2953.LUT_SIZE = 7;
	defparam lut_2953.mask = 128'h77777f7f77777f7f0000153700000000;

	lut_sub lut_2957 ({sk[897], i_5_, i_14_, i_12_, i_11_, x92x, x319x}, x1476x);
	defparam lut_2957.LUT_SIZE = 7;
	defparam lut_2957.mask = 128'h77777f7f77777f7f1111111000000000;

	lut_sub lut_2961 ({sk[898], i_28_, i_29_, x361x, x457x, x388x, x8535x}, x7135x);
	defparam lut_2961.LUT_SIZE = 7;
	defparam lut_2961.mask = 128'h77777f7f77777f7f222f222222222222;

	lut_sub lut_2964 ({sk[899], i_12_, i_11_, x317x, n_n926, x425x, x388x}, x1475x);
	defparam lut_2964.LUT_SIZE = 7;
	defparam lut_2964.mask = 128'h77777f7f77777f7f0007000500070000;

	lut_sub lut_2968 ({sk[900], i_4_, i_1_}, x58x);
	defparam lut_2968.LUT_SIZE = 3;
	defparam lut_2968.mask = 8'h3e;

	lut_sub lut_2971 ({sk[901], i_40_, i_39_, i_34_, i_36_, i_35_, i_38_}, x1469x);
	defparam lut_2971.LUT_SIZE = 7;
	defparam lut_2971.mask = 128'h77777f7f77777f7f0000000000000080;

	lut_sub lut_2973 ({sk[902], i_40_, i_39_, i_38_, i_37_}, x785x);
	defparam lut_2973.LUT_SIZE = 5;
	defparam lut_2973.mask = 32'h00ff080a;

	lut_sub lut_2976 ({sk[903], n_n1055, n_n1047, n_n1048, n_n907, x356x, x785x}, x1467x);
	defparam lut_2976.LUT_SIZE = 7;
	defparam lut_2976.mask = 128'h77777f7f77777f7f000300070003000f;

	lut_sub lut_2980 ({sk[904], i_3_, i_4_, i_1_, i_2_, i_0_, i_32_}, x472x);
	defparam lut_2980.LUT_SIZE = 7;
	defparam lut_2980.mask = 128'h77777f7f77777f7f0000002000000000;

	lut_sub lut_2982 ({sk[905], i_40_, i_14_, i_39_, i_36_, i_38_}, x1463x);
	defparam lut_2982.LUT_SIZE = 6;
	defparam lut_2982.mask = 64'h55ffffff00000400;

	lut_sub lut_2984 ({sk[906], i_40_, i_39_, i_36_, i_38_}, x7148x);
	defparam lut_2984.LUT_SIZE = 5;
	defparam lut_2984.mask = 32'h00ff2000;

	lut_sub lut_2986 ({sk[907], x80x, x7145x, n_n1023, x7147x, x472x, x7148x}, x7152x);
	defparam lut_2986.LUT_SIZE = 7;
	defparam lut_2986.mask = 128'h77777f7f77777f7f0011001100110f1f;

	lut_sub lut_2989 ({sk[908], i_40_, i_39_, i_13_, i_36_, i_38_}, x1071x);
	defparam lut_2989.LUT_SIZE = 6;
	defparam lut_2989.mask = 64'h55ffffff00000800;

	lut_sub lut_2991 ({sk[909], i_39_, i_36_, i_38_, i_37_}, x792x);
	defparam lut_2991.LUT_SIZE = 5;
	defparam lut_2991.mask = 32'h00ff4080;

	lut_sub lut_2994 ({sk[910], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x827x);
	defparam lut_2994.LUT_SIZE = 7;
	defparam lut_2994.mask = 128'h77777f7f77777f7f620080004000a000;

	lut_sub lut_2999 ({sk[911], i_40_, i_39_, i_11_, i_38_, i_37_}, x7078x);
	defparam lut_2999.LUT_SIZE = 6;
	defparam lut_2999.mask = 64'h55ffffff00000008;

	lut_sub lut_3001 ({sk[912], i_6_, i_38_, i_37_, n_n1002, x46x, n_n998}, x1449x);
	defparam lut_3001.LUT_SIZE = 7;
	defparam lut_3001.mask = 128'h77777f7f77777f7f0000000000000311;

	lut_sub lut_3004 ({sk[913], i_12_, n_n990, n_n993, x378x, x76x, x397x}, x7167x);
	defparam lut_3004.LUT_SIZE = 7;
	defparam lut_3004.mask = 128'h77777f7f77777f7f0003000300035557;

	lut_sub lut_3007 ({sk[914], i_5_, i_15_, x422x, x357x, x397x, x7078x}, x7169x);
	defparam lut_3007.LUT_SIZE = 7;
	defparam lut_3007.mask = 128'h77777f7f77777f7f111f111111111111;

	lut_sub lut_3010 ({sk[915], i_6_, x324x, n_n866, n_n884, x336x, x184x}, x8537x);
	defparam lut_3010.LUT_SIZE = 7;
	defparam lut_3010.mask = 128'h77777f7f77777f7fa8a8a8a8a8a8a800;

	lut_sub lut_3017 ({sk[916], i_40_, x1449x, x7167x, x7169x, x8537x}, n_n1675);
	defparam lut_3017.LUT_SIZE = 6;
	defparam lut_3017.mask = 64'h55ffffffbbbbbfff;

	lut_sub lut_3022 ({sk[917], i_40_, i_39_, i_38_, x90x, x51x, x503x}, x802x);
	defparam lut_3022.LUT_SIZE = 7;
	defparam lut_3022.mask = 128'h77777f7f77777f7f550000330f000033;

	lut_sub lut_3026 ({sk[918], x391x, n_n1011, n_n1061, x6797x, x427x, x187x}, x8536x);
	defparam lut_3026.LUT_SIZE = 7;
	defparam lut_3026.mask = 128'h77777f7f77777f7faa80aa80aa800000;

	lut_sub lut_3031 ({sk[919], i_5_, i_13_, i_15_, x7162x, x802x, x8536x}, x7176x);
	defparam lut_3031.LUT_SIZE = 7;
	defparam lut_3031.mask = 128'h77777f7f77777f7fbfafafafafafafaf;

	lut_sub lut_3035 ({sk[920], i_40_, i_39_, i_36_, i_38_, i_37_}, x830x);
	defparam lut_3035.LUT_SIZE = 6;
	defparam lut_3035.mask = 64'h55ffffff80200000;

	lut_sub lut_3038 ({sk[921], i_40_, i_39_, i_36_, i_38_, i_37_}, x829x);
	defparam lut_3038.LUT_SIZE = 6;
	defparam lut_3038.mask = 64'h55ffffff80004000;

	lut_sub lut_3041 ({sk[922], i_22_, x329x, x50x, x87x, x830x, x829x}, x6958x);
	defparam lut_3041.LUT_SIZE = 7;
	defparam lut_3041.mask = 128'h77777f7f77777f7f0005003700000033;

	lut_sub lut_3044 ({sk[923], i_9_, i_39_, i_38_, n_n1047, n_n715, x464x}, x810x);
	defparam lut_3044.LUT_SIZE = 7;
	defparam lut_3044.mask = 128'h77777f7f77777f7f0011001f00110011;

	lut_sub lut_3047 ({sk[924], i_9_, i_5_, i_12_, i_11_, n_n933, n_n927}, x813x);
	defparam lut_3047.LUT_SIZE = 7;
	defparam lut_3047.mask = 128'h77777f7f77777f7f0000000077300000;

	lut_sub lut_3051 ({sk[925], i_9_, i_5_, i_11_, n_n1066, n_n927, x813x}, x812x);
	defparam lut_3051.LUT_SIZE = 7;
	defparam lut_3051.mask = 128'h77777f7f77777f7f0505050507050505;

	lut_sub lut_3054 ({sk[926], i_5_, n_n964, n_n971, n_n977, x404x, x55x}, x817x);
	defparam lut_3054.LUT_SIZE = 7;
	defparam lut_3054.mask = 128'h77777f7f77777f7f000f000f000f777f;

	lut_sub lut_3058 ({sk[927], i_9_, i_32_, i_31_, i_34_, i_33_}, x452x);
	defparam lut_3058.LUT_SIZE = 6;
	defparam lut_3058.mask = 64'h55ffffff00004000;

	lut_sub lut_3060 ({sk[928], i_39_, i_38_, i_37_, n_n1002, x46x, n_n998}, x819x);
	defparam lut_3060.LUT_SIZE = 7;
	defparam lut_3060.mask = 128'h77777f7f77777f7f0003000000000311;

	lut_sub lut_3064 ({sk[929], i_17_, i_15_, i_32_, i_31_, i_34_, i_33_}, x381x);
	defparam lut_3064.LUT_SIZE = 7;
	defparam lut_3064.mask = 128'h77777f7f77777f7f0000400000000000;

	lut_sub lut_3066 ({sk[930], i_7_, i_5_, i_12_, i_11_, i_18_, i_15_}, x1657x);
	defparam lut_3066.LUT_SIZE = 7;
	defparam lut_3066.mask = 128'h77777f7f77777f7f0444000000000000;

	lut_sub lut_3069 ({sk[931], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x605x);
	defparam lut_3069.LUT_SIZE = 7;
	defparam lut_3069.mask = 128'h77777f7f77777f7fb000f000b000d000;

	lut_sub lut_3075 ({sk[932], i_32_, i_34_, i_33_, i_36_, i_35_, i_37_}, x636x);
	defparam lut_3075.LUT_SIZE = 7;
	defparam lut_3075.mask = 128'h77777f7f77777f7f0001008000000000;

	lut_sub lut_3078 ({sk[933], i_40_, i_9_, i_39_, i_13_, i_38_, i_37_}, x659x);
	defparam lut_3078.LUT_SIZE = 7;
	defparam lut_3078.mask = 128'h77777f7f77777f7f000000220c000c22;

	lut_sub lut_3081 ({sk[934], i_30_, i_7_, i_5_, i_28_, i_29_}, x747x);
	defparam lut_3081.LUT_SIZE = 6;
	defparam lut_3081.mask = 64'h55ffffff7000f000;

	lut_sub lut_3085 ({sk[935], i_40_, i_39_, i_36_, i_35_, i_38_, i_37_}, x801x);
	defparam lut_3085.LUT_SIZE = 7;
	defparam lut_3085.mask = 128'h77777f7f77777f7f400080004000a000;

	lut_sub lut_3089 ({sk[936], i_34_, i_36_, i_37_}, x7803x);
	defparam lut_3089.LUT_SIZE = 4;
	defparam lut_3089.mask = 16'h1520;

	lut_sub lut_3091 ({sk[937], i_7_, i_5_, i_12_}, x7796x);
	defparam lut_3091.LUT_SIZE = 4;
	defparam lut_3091.mask = 16'h1580;

	lut_sub lut_3093 ({sk[938], i_40_, i_32_, i_33_, n_n979, n_n975, x315x}, x199x);
	defparam lut_3093.LUT_SIZE = 7;
	defparam lut_3093.mask = 128'h77777f7f77777f7f0000000000010000;

	lut_sub lut_3095 ({sk[939], i_39_, i_38_, i_37_, n_n998, n_n330, n_n700}, x209x);
	defparam lut_3095.LUT_SIZE = 7;
	defparam lut_3095.mask = 128'h77777f7f77777f7f0000000000010000;

	lut_sub lut_3097 ({sk[940], i_36_, i_38_, n_n1014, x69x, x426x, x332x}, x216x);
	defparam lut_3097.LUT_SIZE = 7;
	defparam lut_3097.mask = 128'h77777f7f77777f7f000000000000007f;

	lut_sub lut_3101 ({sk[941], i_5_, i_13_, i_12_}, x7760x);
	defparam lut_3101.LUT_SIZE = 4;
	defparam lut_3101.mask = 16'h1580;

	lut_sub lut_3103 ({sk[942], i_35_, x46x, x323x, x359x, n_n884, x7760x}, x218x);
	defparam lut_3103.LUT_SIZE = 7;
	defparam lut_3103.mask = 128'h77777f7f77777f7f0000073700000000;

	lut_sub lut_3107 ({sk[943], i_3_, i_0_, i_32_, n_n1023, x403x, x58x}, x230x);
	defparam lut_3107.LUT_SIZE = 7;
	defparam lut_3107.mask = 128'h77777f7f77777f7f0000010000000300;

	lut_sub lut_3110 ({sk[944], i_18_, i_21_, i_15_, n_n492, n_n488, x303x}, x275x);
	defparam lut_3110.LUT_SIZE = 7;
	defparam lut_3110.mask = 128'h77777f7f77777f7f0015000000000000;

	lut_sub lut_3113 ({sk[945], i_40_, i_39_, i_38_, i_37_, x513x, x421x}, x295x);
	defparam lut_3113.LUT_SIZE = 7;
	defparam lut_3113.mask = 128'h77777f7f77777f7f0000000000000010;

	lut_sub lut_3115 ({sk[946], i_40_, i_39_, n_n1074, n_n710, n_n1065, x636x}, x311x);
	defparam lut_3115.LUT_SIZE = 7;
	defparam lut_3115.mask = 128'h77777f7f77777f7f0505000000000003;

	lut_sub lut_3118 ({sk[947], i_23_, i_32_, i_33_}, x7694x);
	defparam lut_3118.LUT_SIZE = 4;
	defparam lut_3118.mask = 16'h1540;

	lut_sub lut_3120 ({sk[948], i_5_, i_12_, i_15_, i_32_, i_33_, i_35_}, x7687x);
	defparam lut_3120.LUT_SIZE = 7;
	defparam lut_3120.mask = 128'h77777f7f77777f7f0020000000000000;

	lut_sub lut_3122 ({sk[949], n_n979, n_n853, n_n850, n_n945, n_n848, n_n866}, x466x);
	defparam lut_3122.LUT_SIZE = 7;
	defparam lut_3122.mask = 128'h77777f7f77777f7f0000000000010101;

	lut_sub lut_3125 ({sk[950], i_40_, i_39_, i_38_, x35x, n_n848, x340x}, x477x);
	defparam lut_3125.LUT_SIZE = 7;
	defparam lut_3125.mask = 128'h77777f7f77777f7f0000000000000100;

	lut_sub lut_3127 ({sk[951], i_24_, i_32_, x82x, n_n528, x87x, n_n1023}, x519x);
	defparam lut_3127.LUT_SIZE = 7;
	defparam lut_3127.mask = 128'h77777f7f77777f7f0000000001050000;

	lut_sub lut_3130 ({sk[952], i_32_, i_31_, n_n462, n_n1066, x102x}, x858x);
	defparam lut_3130.LUT_SIZE = 6;
	defparam lut_3130.mask = 64'h55ffffff01000000;

	lut_sub lut_3132 ({sk[953], i_7_, i_4_, i_1_, i_0_, n_n1074}, x8555x);
	defparam lut_3132.LUT_SIZE = 6;
	defparam lut_3132.mask = 64'h55ffffffeeefffff;

	lut_sub lut_3137 ({sk[954], i_40_, i_35_, i_38_, i_37_, x302x, x8555x}, x891x);
	defparam lut_3137.LUT_SIZE = 7;
	defparam lut_3137.mask = 128'h77777f7f77777f7f00000b0000000000;

	lut_sub lut_3140 ({sk[955], i_4_, i_1_, i_0_, x302x, x79x, x402x}, x892x);
	defparam lut_3140.LUT_SIZE = 7;
	defparam lut_3140.mask = 128'h77777f7f77777f7f0505051505150515;

	lut_sub lut_3144 ({sk[956], i_7_, i_5_, i_12_, i_11_, i_32_, i_31_}, x7609x);
	defparam lut_3144.LUT_SIZE = 7;
	defparam lut_3144.mask = 128'h77777f7f77777f7f8000000000000000;

	lut_sub lut_3146 ({sk[957], n_n330, x325x, n_n989, x445x, n_n976, x7609x}, x912x);
	defparam lut_3146.LUT_SIZE = 7;
	defparam lut_3146.mask = 128'h77777f7f77777f7f0000111100031113;

	lut_sub lut_3149 ({sk[958], i_12_, i_11_, i_15_, x47x, x93x, n_n469}, x913x);
	defparam lut_3149.LUT_SIZE = 7;
	defparam lut_3149.mask = 128'h77777f7f77777f7f0101010101010100;

	lut_sub lut_3153 ({sk[959], i_40_, i_36_, i_35_, i_38_, i_37_, x429x}, x926x);
	defparam lut_3153.LUT_SIZE = 7;
	defparam lut_3153.mask = 128'h77777f7f77777f7f0010001000000500;

	lut_sub lut_3156 ({sk[960], i_34_, n_n1021, x81x, n_n1048, x398x, x747x}, x927x);
	defparam lut_3156.LUT_SIZE = 7;
	defparam lut_3156.mask = 128'h77777f7f77777f7f0000333700003333;

	lut_sub lut_3159 ({sk[961], i_14_, n_n853, n_n775, n_n1048, x78x, x327x}, x942x);
	defparam lut_3159.LUT_SIZE = 7;
	defparam lut_3159.mask = 128'h77777f7f77777f7f0000010300000000;

	lut_sub lut_3162 ({sk[962], i_18_, i_19_, i_37_, n_n1011, x6977x, x486x}, x943x);
	defparam lut_3162.LUT_SIZE = 7;
	defparam lut_3162.mask = 128'h77777f7f77777f7f0001000000000000;

	lut_sub lut_3164 ({sk[963], x82x, n_n775, n_n1048, x87x, x37x, x327x}, x944x);
	defparam lut_3164.LUT_SIZE = 7;
	defparam lut_3164.mask = 128'h77777f7f77777f7f0004000c004400cc;

	lut_sub lut_3169 ({sk[964], i_40_, n_n761, n_n833, n_n764, n_n836, n_n765}, x962x);
	defparam lut_3169.LUT_SIZE = 7;
	defparam lut_3169.mask = 128'h77777f7f77777f7f135f33ff005f00ff;

	lut_sub lut_3176 ({sk[965], i_7_, i_25_, i_26_, i_32_, n_n1023, n_n693}, x986x);
	defparam lut_3176.LUT_SIZE = 7;
	defparam lut_3176.mask = 128'h77777f7f77777f7f1000101000000000;

	lut_sub lut_3179 ({sk[966], i_5_, n_n968, x480x, x120x, x86x, x78x}, x997x);
	defparam lut_3179.LUT_SIZE = 7;
	defparam lut_3179.mask = 128'h77777f7f77777f7f0000000700000000;

	lut_sub lut_3182 ({sk[967], i_5_, i_12_, i_11_, i_15_, x52x, x7134x}, x998x);
	defparam lut_3182.LUT_SIZE = 7;
	defparam lut_3182.mask = 128'h77777f7f77777f7f0001010100000000;

	lut_sub lut_3185 ({sk[968], i_9_, i_7_, i_17_, i_16_, i_38_, x424x}, x1049x);
	defparam lut_3185.LUT_SIZE = 7;
	defparam lut_3185.mask = 128'h77777f7f77777f7f4440000040000000;

	lut_sub lut_3189 ({sk[969], i_7_, i_15_, x45x, x50x, x101x, x357x}, x1050x);
	defparam lut_3189.LUT_SIZE = 7;
	defparam lut_3189.mask = 128'h77777f7f77777f7f0357000000000000;

	lut_sub lut_3192 ({sk[970], i_40_, i_39_, i_24_, i_38_, x51x, x365x}, x1121x);
	defparam lut_3192.LUT_SIZE = 7;
	defparam lut_3192.mask = 128'h77777f7f77777f7f0010000100000000;

	lut_sub lut_3195 ({sk[971], i_4_, i_0_, i_32_, i_36_, n_n1023, x403x}, x1155x);
	defparam lut_3195.LUT_SIZE = 7;
	defparam lut_3195.mask = 128'h77777f7f77777f7f0000010000000000;

	lut_sub lut_3197 ({sk[972], i_21_, i_22_, x46x, n_n1001, x338x, x360x}, x1187x);
	defparam lut_3197.LUT_SIZE = 7;
	defparam lut_3197.mask = 128'h77777f7f77777f7f0007000700070000;

	lut_sub lut_3202 ({sk[973], i_4_, i_1_, x95x, x429x, x350x, x302x}, x1213x);
	defparam lut_3202.LUT_SIZE = 7;
	defparam lut_3202.mask = 128'h77777f7f77777f7f007f007f007f005f;

	lut_sub lut_3207 ({sk[974], i_7_, i_32_, i_33_, n_n969, n_n971, x7334x}, x1254x);
	defparam lut_3207.LUT_SIZE = 7;
	defparam lut_3207.mask = 128'h77777f7f77777f7f0057000000000000;

	lut_sub lut_3210 ({sk[975], i_40_, i_39_, i_35_, i_38_, i_37_, x411x}, x1273x);
	defparam lut_3210.LUT_SIZE = 7;
	defparam lut_3210.mask = 128'h77777f7f77777f7f0010000000000000;

	lut_sub lut_3212 ({sk[976], i_14_, i_17_, i_16_, n_n560, x327x, x41x}, x8549x);
	defparam lut_3212.LUT_SIZE = 7;
	defparam lut_3212.mask = 128'h77777f7f77777f7f00000000002a2a2a;

	lut_sub lut_3217 ({sk[977], i_40_, i_30_, i_39_, i_38_, n_n1047, x494x}, x8528x);
	defparam lut_3217.LUT_SIZE = 7;
	defparam lut_3217.mask = 128'h77777f7f77777f7ffffffffffeffffff;

	lut_sub lut_3232 ({sk[978], i_35_, i_38_, i_37_, n_n1074, n_n710, x89x}, x1333x);
	defparam lut_3232.LUT_SIZE = 7;
	defparam lut_3232.mask = 128'h77777f7f77777f7f1111111111111113;

	lut_sub lut_3235 ({sk[979], i_3_, i_4_, i_1_, i_38_, i_37_, x77x}, x1341x);
	defparam lut_3235.LUT_SIZE = 7;
	defparam lut_3235.mask = 128'h77777f7f77777f7f0010101010101010;

	lut_sub lut_3239 ({sk[980], i_40_, i_32_, i_34_, i_33_, i_36_, i_35_}, x1361x);
	defparam lut_3239.LUT_SIZE = 7;
	defparam lut_3239.mask = 128'h77777f7f77777f7f0200000000000000;

	lut_sub lut_3241 ({sk[981], i_14_, i_12_, x317x, n_n926, x425x, x1463x}, x1460x);
	defparam lut_3241.LUT_SIZE = 7;
	defparam lut_3241.mask = 128'h77777f7f77777f7f0013001300130011;

	lut_sub lut_3245 ({sk[982], i_5_, i_14_, i_12_, i_11_, n_n926, x319x}, x1461x);
	defparam lut_3245.LUT_SIZE = 7;
	defparam lut_3245.mask = 128'h77777f7f77777f7f1111111000000000;

	lut_sub lut_3249 ({sk[983], i_36_, n_n1067, x100x, n_n1023, n_n1057, x393x}, x1466x);
	defparam lut_3249.LUT_SIZE = 7;
	defparam lut_3249.mask = 128'h77777f7f77777f7f0000555500005557;

	lut_sub lut_3252 ({sk[984], i_40_, i_39_, i_34_, i_36_, i_38_, i_37_}, x1514x);
	defparam lut_3252.LUT_SIZE = 7;
	defparam lut_3252.mask = 128'h77777f7f77777f7f0000000001000000;

	lut_sub lut_3254 ({sk[985], i_40_, i_39_, i_38_, n_n979, n_n980, n_n1012}, x1523x);
	defparam lut_3254.LUT_SIZE = 7;
	defparam lut_3254.mask = 128'h77777f7f77777f7f0000000003001100;

	lut_sub lut_3257 ({sk[986], n_n1006, n_n983, x7090x, n_n977, n_n1023, n_n1065}, x1524x);
	defparam lut_3257.LUT_SIZE = 7;
	defparam lut_3257.mask = 128'h77777f7f77777f7f0000000011ff1fff;

	lut_sub lut_3261 ({sk[987], i_39_, i_15_, i_36_, i_35_, i_37_, x452x}, x1539x);
	defparam lut_3261.LUT_SIZE = 7;
	defparam lut_3261.mask = 128'h77777f7f77777f7f0000000040000000;

	lut_sub lut_3263 ({sk[988], i_40_, i_3_, i_39_, i_4_, n_n1061, n_n1065}, x8548x);
	defparam lut_3263.LUT_SIZE = 7;
	defparam lut_3263.mask = 128'h77777f7f77777f7fffcfffffafcfffff;

	lut_sub lut_3283 ({sk[989], i_14_, i_17_, i_16_, i_31_, x46x, n_n775}, x1566x);
	defparam lut_3283.LUT_SIZE = 7;
	defparam lut_3283.mask = 128'h77777f7f77777f7f0000001000000000;

	lut_sub lut_3285 ({sk[990], i_9_, i_14_, i_12_, i_11_, i_17_, i_16_}, x7051x);
	defparam lut_3285.LUT_SIZE = 7;
	defparam lut_3285.mask = 128'h77777f7f77777f7f1110111033333130;

	lut_sub lut_3290 ({sk[991], i_5_, i_14_, i_12_, i_11_, i_15_, x91x}, x1583x);
	defparam lut_3290.LUT_SIZE = 7;
	defparam lut_3290.mask = 128'h77777f7f77777f7f0000000055555554;

	lut_sub lut_3295 ({sk[992], i_17_, i_16_, x82x, n_n775, n_n1048, x87x}, x1717x);
	defparam lut_3295.LUT_SIZE = 7;
	defparam lut_3295.mask = 128'h77777f7f77777f7f0103000000000000;

	lut_sub lut_3298 ({sk[993], i_12_, i_18_, i_24_, i_22_, x35x, n_n793}, x8552x);
	defparam lut_3298.LUT_SIZE = 7;
	defparam lut_3298.mask = 128'h77777f7f77777f7ffffcfffffff8fffa;

	lut_sub lut_3315 ({sk[994], n_n979, n_n945, x400x, n_n528, n_n902, x36x}, x6718x);
	defparam lut_3315.LUT_SIZE = 7;
	defparam lut_3315.mask = 128'h77777f7f77777f7f0033003300330537;

	lut_sub lut_3318 ({sk[995], n_n979, n_n973, n_n1012, n_n866, x399x, x356x}, x6746x);
	defparam lut_3318.LUT_SIZE = 7;
	defparam lut_3318.mask = 128'h77777f7f77777f7f1111113313131333;

	lut_sub lut_3322 ({sk[996], i_15_, n_n955, n_n1159, x66x, x90x, x537x}, x8546x);
	defparam lut_3322.LUT_SIZE = 7;
	defparam lut_3322.mask = 128'h77777f7f77777f7ffc00fc00fc00a800;

	lut_sub lut_3329 ({sk[997], i_40_, i_39_, i_38_, n_n1074, n_n1061, n_n970}, x6803x);
	defparam lut_3329.LUT_SIZE = 7;
	defparam lut_3329.mask = 128'h77777f7f77777f7f0000050007030500;

	lut_sub lut_3333 ({sk[998], i_25_, i_26_, x530x, x340x, n_n799, x187x}, x8545x);
	defparam lut_3333.LUT_SIZE = 7;
	defparam lut_3333.mask = 128'h77777f7f77777f7fa8a8a800a800a800;

	lut_sub lut_3338 ({sk[999], i_40_, i_39_, i_38_, x90x, x391x, x89x}, x8551x);
	defparam lut_3338.LUT_SIZE = 7;
	defparam lut_3338.mask = 128'h77777f7f77777f7ff0aaffccfffffff0;

	lut_sub lut_3350 ({sk[1000], i_40_, i_13_, x47x, n_n926, n_n1009, x387x}, x6875x);
	defparam lut_3350.LUT_SIZE = 7;
	defparam lut_3350.mask = 128'h77777f7f77777f7f0000001500000005;

	lut_sub lut_3353 ({sk[1001], x366x, n_n775, n_n1048, x76x, x6856x, x6834x}, x6909x);
	defparam lut_3353.LUT_SIZE = 7;
	defparam lut_3353.mask = 128'h77777f7f77777f7f0000003305050537;

	lut_sub lut_3356 ({sk[1002], i_17_, i_16_, n_n775, n_n1048, x1787x, x367x}, x6910x);
	defparam lut_3356.LUT_SIZE = 7;
	defparam lut_3356.mask = 128'h77777f7f77777f7f0105000501050000;

	lut_sub lut_3360 ({sk[1003], i_40_, i_39_, n_n985, x329x, n_n1983, x80x}, x6956x);
	defparam lut_3360.LUT_SIZE = 7;
	defparam lut_3360.mask = 128'h77777f7f77777f7f3333333333333337;

	lut_sub lut_3363 ({sk[1004], x93x, x50x, x6955x, x87x, x367x, x6859x}, x6957x);
	defparam lut_3363.LUT_SIZE = 7;
	defparam lut_3363.mask = 128'h77777f7f77777f7f0000000f1111111f;

	lut_sub lut_3366 ({sk[1005], i_40_, i_39_, i_38_, i_37_, n_n861, n_n998}, x7020x);
	defparam lut_3366.LUT_SIZE = 7;
	defparam lut_3366.mask = 128'h77777f7f77777f7f0010000000111000;

	lut_sub lut_3370 ({sk[1006], i_23_, i_32_, x329x, x323x, x87x, n_n1023}, x7034x);
	defparam lut_3370.LUT_SIZE = 7;
	defparam lut_3370.mask = 128'h77777f7f77777f7f0105000000050000;

	lut_sub lut_3373 ({sk[1007], n_n985, n_n1064, n_n760, n_n833, n_n764, x101x}, x8558x);
	defparam lut_3373.LUT_SIZE = 7;
	defparam lut_3373.mask = 128'h77777f7f77777f7ffca8fca8fca8fc00;

	lut_sub lut_3380 ({sk[1008], i_40_, i_39_, i_36_, i_38_, x389x, x387x}, x7075x);
	defparam lut_3380.LUT_SIZE = 7;
	defparam lut_3380.mask = 128'h77777f7f77777f7f3030000050005000;

	lut_sub lut_3383 ({sk[1009], i_40_, i_39_, i_38_, n_n1074, n_n968, x340x}, x7076x);
	defparam lut_3383.LUT_SIZE = 7;
	defparam lut_3383.mask = 128'h77777f7f77777f7f0057000000000300;

	lut_sub lut_3387 ({sk[1010], n_n926, n_n989, n_n983, x387x, x445x, x1523x}, x7092x);
	defparam lut_3387.LUT_SIZE = 7;
	defparam lut_3387.mask = 128'h77777f7f77777f7f555555775f5f5f7f;

	lut_sub lut_3391 ({sk[1011], i_40_, i_14_, i_36_, x317x, n_n926, n_n960}, x8535x);
	defparam lut_3391.LUT_SIZE = 7;
	defparam lut_3391.mask = 128'h77777f7f77777f7ffcfcfffff8fcffff;

	lut_sub lut_3405 ({sk[1012], n_n979, n_n969, n_n1001, n_n888, x399x, x1469x}, x7143x);
	defparam lut_3405.LUT_SIZE = 7;
	defparam lut_3405.mask = 128'h77777f7f77777f7f1111131311331333;

	lut_sub lut_3409 ({sk[1013], i_40_, i_5_, i_38_, x93x, x61x, x140x}, x7174x);
	defparam lut_3409.LUT_SIZE = 7;
	defparam lut_3409.mask = 128'h77777f7f77777f7f555555555d555555;

	lut_sub lut_3412 ({sk[1014], x317x, x378x, x76x, x521x, x801x, x7174x}, x7175x);
	defparam lut_3412.LUT_SIZE = 7;
	defparam lut_3412.mask = 128'h77777f7f77777f7f55555577555f557f;

	lut_sub lut_3416 ({sk[1015], i_12_, i_11_, i_15_, i_37_, x317x, x490x}, x8534x);
	defparam lut_3416.LUT_SIZE = 7;
	defparam lut_3416.mask = 128'h77777f7f77777f7fefefefefefefefff;

	lut_sub lut_3429 ({sk[1016], i_40_, n_n1055, n_n977, n_n1048, n_n902, x8534x}, x7183x);
	defparam lut_3429.LUT_SIZE = 7;
	defparam lut_3429.mask = 128'h77777f7f77777f7f000a333b000a000a;

	lut_sub lut_3432 ({sk[1017], i_40_, i_39_, i_38_, i_37_, x354x, x392x}, x7219x);
	defparam lut_3432.LUT_SIZE = 7;
	defparam lut_3432.mask = 128'h77777f7f77777f7f7557555555550000;

	lut_sub lut_3437 ({sk[1018], x330x, x335x, n_n685, x7212x, x251x, x7219x}, x7222x);
	defparam lut_3437.LUT_SIZE = 7;
	defparam lut_3437.mask = 128'h77777f7f77777f7f777777ff7f7f7fff;

	lut_sub lut_3442 ({sk[1019], i_9_, i_5_, i_32_, x49x, x110x, x750x}, x8532x);
	defparam lut_3442.LUT_SIZE = 7;
	defparam lut_3442.mask = 128'h77777f7f77777f7ffff0f8f0fff0faf0;

	lut_sub lut_3447 ({sk[1020], i_32_, i_33_, x51x, n_n960, n_n1073, x41x}, x7243x);
	defparam lut_3447.LUT_SIZE = 7;
	defparam lut_3447.mask = 128'h77777f7f77777f7f000f010f000f000f;

	lut_sub lut_3450 ({sk[1021], i_39_, i_38_, n_n1074, n_n971, n_n1047, n_n700}, x7244x);
	defparam lut_3450.LUT_SIZE = 7;
	defparam lut_3450.mask = 128'h77777f7f77777f7f0000000f11110000;

	lut_sub lut_3453 ({sk[1022], i_5_, i_34_, i_36_, i_35_, i_38_, x46x}, x7266x);
	defparam lut_3453.LUT_SIZE = 7;
	defparam lut_3453.mask = 128'h77777f7f77777f7f0000000050100000;

	lut_sub lut_3456 ({sk[1023], i_7_, i_33_, n_n1014, n_n966, n_n862, x339x}, x7267x);
	defparam lut_3456.LUT_SIZE = 7;
	defparam lut_3456.mask = 128'h77777f7f77777f7f575557555755ffff;

	lut_sub lut_3460 ({sk[1024], i_38_, x90x, x391x, n_n1021, x89x, x413x}, x8530x);
	defparam lut_3460.LUT_SIZE = 7;
	defparam lut_3460.mask = 128'h77777f7f77777f7faa000a0088880808;

	lut_sub lut_3467 ({sk[1025], i_31_, n_n1008, x47x, n_n1066, n_n1052, n_n582}, x8527x);
	defparam lut_3467.LUT_SIZE = 7;
	defparam lut_3467.mask = 128'h77777f7f77777f7ffffffff8ffffffff;

	lut_sub lut_3482 ({sk[1026], i_40_, i_31_, i_34_, i_33_}, x7314x);
	defparam lut_3482.LUT_SIZE = 5;
	defparam lut_3482.mask = 32'h00ff4000;

	lut_sub lut_3484 ({sk[1027], i_38_, i_37_, x88x, n_n1021, n_n979, x328x}, x7335x);
	defparam lut_3484.LUT_SIZE = 7;
	defparam lut_3484.mask = 128'h77777f7f77777f7f0000053700000505;

	lut_sub lut_3487 ({sk[1028], i_39_, i_38_, i_37_, n_n979, n_n861, x177x}, x7336x);
	defparam lut_3487.LUT_SIZE = 7;
	defparam lut_3487.mask = 128'h77777f7f77777f7f5555555755555555;

	lut_sub lut_3490 ({sk[1029], i_39_, i_32_, i_38_, n_n861, n_n998, x49x}, x7343x);
	defparam lut_3490.LUT_SIZE = 7;
	defparam lut_3490.mask = 128'h77777f7f77777f7f0003555700005555;

	lut_sub lut_3493 ({sk[1030], n_n979, x335x, n_n469, x396x, x364x, x7347x}, x8565x);
	defparam lut_3493.LUT_SIZE = 7;
	defparam lut_3493.mask = 128'h77777f7f77777f7ffffff0f0ffeef0e0;

	lut_sub lut_3502 ({sk[1031], i_40_, i_39_, n_n862, x76x, x6834x, x6862x}, x7377x);
	defparam lut_3502.LUT_SIZE = 7;
	defparam lut_3502.mask = 128'h77777f7f77777f7f0000000000070000;

	lut_sub lut_3505 ({sk[1032], i_22_, x82x, x50x, n_n833, x245x, x87x}, x8557x);
	defparam lut_3505.LUT_SIZE = 7;
	defparam lut_3505.mask = 128'h77777f7f77777f7fccc8ccc0cccccccc;

	lut_sub lut_3510 ({sk[1033], i_24_, i_32_, i_33_, i_38_, n_n1064, x65x}, x8574x);
	defparam lut_3510.LUT_SIZE = 7;
	defparam lut_3510.mask = 128'h77777f7f77777f7fff8affffffffffff;

	lut_sub lut_3525 ({sk[1034], i_28_, i_29_, x361x, x406x, x338x, x8574x}, x7410x);
	defparam lut_3525.LUT_SIZE = 7;
	defparam lut_3525.mask = 128'h77777f7f77777f7f22222222222f2222;

	lut_sub lut_3528 ({sk[1035], i_39_, i_37_, n_n964, n_n488, x401x, x352x}, x8573x);
	defparam lut_3528.LUT_SIZE = 7;
	defparam lut_3528.mask = 128'h77777f7f77777f7ffefefefefefafefe;

	lut_sub lut_3542 ({sk[1036], i_36_, x502x, n_n799, x403x, x680x, x1155x}, x8523x);
	defparam lut_3542.LUT_SIZE = 7;
	defparam lut_3542.mask = 128'h77777f7f77777f7faaaaaa00a8a8a800;

	lut_sub lut_3549 ({sk[1037], i_7_, i_4_, i_33_, x384x, x69x, x394x}, x8524x);
	defparam lut_3549.LUT_SIZE = 7;
	defparam lut_3549.mask = 128'h77777f7f77777f7feeeee0e0ee00e000;

	lut_sub lut_3558 ({sk[1038], n_n1983, n_n1927, n_n1980, x1121x}, x7462x);
	defparam lut_3558.LUT_SIZE = 5;
	defparam lut_3558.mask = 32'h00ff7fff;

	lut_sub lut_3563 ({sk[1039], i_36_, x390x, x182x, x301x, x7468x, x659x}, x8521x);
	defparam lut_3563.LUT_SIZE = 7;
	defparam lut_3563.mask = 128'h77777f7f77777f7ff0008000f000c000;

	lut_sub lut_3567 ({sk[1040], i_7_, n_n1074, n_n560, x61x, x303x, x233x}, x8567x);
	defparam lut_3567.LUT_SIZE = 7;
	defparam lut_3567.mask = 128'h77777f7f77777f7f8f8f8f0fffffffff;

	lut_sub lut_3580 ({sk[1041], i_37_, n_n1021, n_n861, x358x, n_n799, x624x}, x7552x);
	defparam lut_3580.LUT_SIZE = 7;
	defparam lut_3580.mask = 128'h77777f7f77777f7f00110f1f00110011;

	lut_sub lut_3583 ({sk[1042], i_39_, i_38_, i_37_, x88x, n_n979, x358x}, x7553x);
	defparam lut_3583.LUT_SIZE = 7;
	defparam lut_3583.mask = 128'h77777f7f77777f7f0003000055030000;

	lut_sub lut_3586 ({sk[1043], i_7_, i_5_, i_29_, x181x, n_n462, x361x}, x7596x);
	defparam lut_3586.LUT_SIZE = 7;
	defparam lut_3586.mask = 128'h77777f7f77777f7f1f0f0f0f0f0f0f0f;

	lut_sub lut_3589 ({sk[1044], i_36_, n_n330, x387x, x68x, n_n287, x124x}, x7597x);
	defparam lut_3589.LUT_SIZE = 7;
	defparam lut_3589.mask = 128'h77777f7f77777f7f1111111f11111111;

	lut_sub lut_3592 ({sk[1045], i_15_, x47x, n_n973, n_n1048, n_n1073, x926x}, x7604x);
	defparam lut_3592.LUT_SIZE = 7;
	defparam lut_3592.mask = 128'h77777f7f77777f7f5555555755555555;

	lut_sub lut_3595 ({sk[1046], x94x, n_n330, n_n926, n_n975, x387x, x97x}, x7611x);
	defparam lut_3595.LUT_SIZE = 7;
	defparam lut_3595.mask = 128'h77777f7f77777f7f0000003305050537;

	lut_sub lut_3598 ({sk[1047], n_n837, n_n834, n_n836, x408x, x76x, x103x}, x8518x);
	defparam lut_3598.LUT_SIZE = 7;
	defparam lut_3598.mask = 128'h77777f7f77777f7ffefefe00fe00fe00;

	lut_sub lut_3605 ({sk[1048], i_7_, i_39_, i_38_, i_37_, x46x, n_n991}, x8568x);
	defparam lut_3605.LUT_SIZE = 7;
	defparam lut_3605.mask = 128'h77777f7f77777f7ffeeffffeffffffff;

	lut_sub lut_3631 ({sk[1049], i_2_, i_0_, n_n1021, x313x, x438x, x493x}, x7634x);
	defparam lut_3631.LUT_SIZE = 7;
	defparam lut_3631.mask = 128'h77777f7f77777f7f0000000533333337;

	lut_sub lut_3634 ({sk[1050], i_40_, i_39_, i_15_, i_38_, i_37_, x47x}, x8564x);
	defparam lut_3634.LUT_SIZE = 7;
	defparam lut_3634.mask = 128'h77777f7f77777f7fffffffffefffbfff;

	lut_sub lut_3651 ({sk[1051], i_13_, x47x, x93x, n_n926, x387x, x8564x}, x7662x);
	defparam lut_3651.LUT_SIZE = 7;
	defparam lut_3651.mask = 128'h77777f7f77777f7f00aa00aa00aa03ab;

	lut_sub lut_3654 ({sk[1052], i_40_, i_13_, i_32_, n_n833, n_n975, n_n1023}, x8572x);
	defparam lut_3654.LUT_SIZE = 7;
	defparam lut_3654.mask = 128'h77777f7f77777f7feafffffffaffffff;

	lut_sub lut_3669 ({sk[1053], x358x, n_n883, n_n462, x361x, n_n710, x494x}, x7672x);
	defparam lut_3669.LUT_SIZE = 7;
	defparam lut_3669.mask = 128'h77777f7f77777f7f0005000500053337;

	lut_sub lut_3672 ({sk[1054], i_39_, i_16_, i_15_, x91x, n_n488, x154x}, x7702x);
	defparam lut_3672.LUT_SIZE = 7;
	defparam lut_3672.mask = 128'h77777f7f77777f7f5555555555575555;

	lut_sub lut_3675 ({sk[1055], i_38_, n_n964, n_n775, x460x, x427x, x635x}, x7703x);
	defparam lut_3675.LUT_SIZE = 7;
	defparam lut_3675.mask = 128'h77777f7f77777f7f000f000f000f111f;

	lut_sub lut_3678 ({sk[1056], i_14_, i_39_, i_17_, i_15_, i_36_, i_38_}, x8570x);
	defparam lut_3678.LUT_SIZE = 7;
	defparam lut_3678.mask = 128'h77777f7f77777f7ffffffbfffffffbfb;

	lut_sub lut_3693 ({sk[1057], i_15_, x92x, x517x, x110x, x331x, x7725x}, x7729x);
	defparam lut_3693.LUT_SIZE = 7;
	defparam lut_3693.mask = 128'h77777f7f77777f7f0033003300335073;

	lut_sub lut_3696 ({sk[1058], i_40_, i_39_, x81x, n_n1023, n_n458, x413x}, x7746x);
	defparam lut_3696.LUT_SIZE = 7;
	defparam lut_3696.mask = 128'h77777f7f77777f7f0003555700000000;

	lut_sub lut_3699 ({sk[1059], i_9_, i_5_, x391x, x45x, n_n997, n_n977}, x7751x);
	defparam lut_3699.LUT_SIZE = 7;
	defparam lut_3699.mask = 128'h77777f7f77777f7f0357005500550055;

	lut_sub lut_3702 ({sk[1060], i_40_, i_39_, i_38_, n_n1074, n_n864, x340x}, x7752x);
	defparam lut_3702.LUT_SIZE = 7;
	defparam lut_3702.mask = 128'h77777f7f77777f7f0000000055030000;

	lut_sub lut_3705 ({sk[1061], i_25_, i_1_, i_37_, x324x, n_n1011, x77x}, x7753x);
	defparam lut_3705.LUT_SIZE = 7;
	defparam lut_3705.mask = 128'h77777f7f77777f7f0300031100000011;

	lut_sub lut_3708 ({sk[1062], x218x, x230x, x7751x, x7752x, x7753x}, x7762x);
	defparam lut_3708.LUT_SIZE = 6;
	defparam lut_3708.mask = 64'h55ffffff7fffffff;

	lut_sub lut_3714 ({sk[1063], i_40_, x45x, x355x, x202x, x406x, x683x}, x8513x);
	defparam lut_3714.LUT_SIZE = 7;
	defparam lut_3714.mask = 128'h77777f7f77777f7ffffffcfcffaafca8;

	lut_sub lut_3724 ({sk[1064], i_7_, i_5_, i_13_, n_n866, n_n700, x65x}, x8556x);
	defparam lut_3724.LUT_SIZE = 7;
	defparam lut_3724.mask = 128'h77777f7f77777f7fffecffffffffffff;


endmodule