module apex2_o (input i_0_, input i_1_, input i_2_, input i_3_, input i_4_, input i_5_, input i_6_, input i_7_, input i_8_, input i_9_, input i_10_, input i_11_, input i_12_, input i_13_, input i_14_, input i_15_, input i_16_, input i_17_, input i_18_, input i_19_, input i_20_, input i_21_, input i_22_, input i_23_, input i_24_, input i_25_, input i_26_, input i_27_, input i_28_, input i_29_, input i_30_, input i_31_, input i_32_, input i_33_, input i_34_, input i_35_, input i_36_, input i_37_, input i_38_, output o_0_, output o_1_, output o_2_);



	wire n1, n2, n3, n5, n8, n1248, n1249, n1250, n753, n433, n245;
	wire n479, n880, n1025, n670, n669, n874, n885, n1035, n216, n608, n662;
	wire n1215, n217, n939, n942, n944, n947, n950, n1033, n1253, n163, n10;
	wire n350, n11, n1213, n9, n15, n1030, n13, n19, n60, n59, n17;
	wire n24, n23, n22, n67, n66, n26, n30, n31, n29, n33, n70;
	wire n32, n35, n966, n769, n38, n256, n39, n97, n40, n36, n44;
	wire n147, n1000, n41, n48, n45, n324, n394, n800, n52, n968, n50;
	wire n121, n49, n90, n135, n56, n290, n402, n53, n990, n371, n84;
	wire n57, n964, n64, n374, n965, n63, n61, n985, n81, n65, n69;
	wire n986, n68, n977, n72, n73, n74, n71, n75, n78, n989, n82;
	wire n299, n80, n91, n322, n87, n100, n88, n963, n86, n85, n89;
	wire n983, n528, n93, n991, n94, n92, n595, n96, n229, n98, n95;
	wire n970, n101, n99, n104, n102, n1258, n107, n105, n1001, n1117, n112;
	wire n110, n1116, n111, n109, n1118, n1121, n1123, n113, n1126, n1129, n1132;
	wire n117, n162, n313, n125, n195, n306, n994, n126, n988, n124, n122;
	wire n179, n129, n288, n130, n138, n131, n127, n133, n134, n132, n139;
	wire n136, n311, n140, n144, n145, n143, n962, n148, n146, n150, n151;
	wire n149, n152, n414, n155, n326, n159, n1115, n160, n157, n161, n367;
	wire n167, n170, n165, n308, n166, n164, n168, n304, n171, n972, n175;
	wire n206, n176, n685, n174, n173, n180, n177, n987, n183, n184, n182;
	wire n181, n185, n188, n189, n190, n429, n186, n193, n234, n192, n191;
	wire n832, n197, n196, n194, n199, n200, n198, n648, n203, n241, n376;
	wire n204, n201, n205, n253, n211, n207, n957, n213, n960, n215, n734;
	wire n363, n212, n681, n954, n219, n673, n222, n221, n224, n225, n227;
	wire n226, n232, n230, n995, n236, n233, n356, n239, n724, n238, n237;
	wire n240, n974, n243, n242, n246, n244, n1012, n248, n249, n247, n250;
	wire n1097, n252, n255, n258, n261, n260, n263, n266, n265, n264, n268;
	wire n267, n269, n272, n273, n274, n282, n279, n1088, n278, n283, n284;
	wire n287, n289, n293, n1057, n296, n300, n301, n307, n305, n309, n315;
	wire n314, n1081, n317, n319, n320, n323, n325, n996, n328, n331, n349;
	wire n1065, n335, n1066, n336, n334, n332, n337, n716, n341, n340, n339;
	wire n342, n978, n345, n346, n347, n344, n348, n1062, n352, n1063, n355;
	wire n1067, n1069, n358, n362, n833, n364, n361, n365, n368, n961, n372;
	wire n373, n370, n375, n377, n1045, n1046, n378, n382, n1047, n1048, n1049;
	wire n1051, n385, n1053, n1055, n1058, n390, n395, n397, n399, n404, n403;
	wire n407, n406, n1089, n1091, n1093, n408, n413, n412, n1263, n415, n1102;
	wire n418, n997, n1106, n421, n1108, n425, n1113, n428, n531, n436, n1141;
	wire n969, n437, n1139, n438, n1146, n439, n1143, n440, n1149, n1152, n1153;
	wire n1157, n1159, n1160, n441, n443, n649, n444, n446, n442, n543, n664;
	wire n449, n448, n447, n451, n450, n453, n1020, n455, n735, n454, n452;
	wire n1015, n522, n501, n459, n622, n457, n1114, n458, n456, n494, n992;
	wire n462, n1005, n461, n460, n467, n629, n1194, n463, n639, n1009, n587;
	wire n471, n469, n746, n470, n468, n474, n692, n473, n953, n688, n477;
	wire n763, n482, n481, n480, n572, n485, n483, n1027, n487, n884, n561;
	wire n1023, n488, n489, n1196, n684, n490, n486, n495, n1011, n491, n497;
	wire n498, n496, n500, n503, n505, n502, n609, n620, n506, n1003, n512;
	wire n513, n511, n1169, n1013, n516, n515, n514, n640, n519, n518, n517;
	wire n520, n521, n1192, n526, n524, n523, n1007, n527, n525, n1190, n529;
	wire n1014, n556, n534, n533, n539, n535, n704, n1193, n540, n1163, n984;
	wire n545, n544, n547, n548, n546, n550, n549, n554, n552, n557, n558;
	wire n559, n555, n607, n562, n717, n560, n1187, n563, n1188, n569, n567;
	wire n841, n573, n570, n586, n576, n1010, n575, n574, n578, n631, n1016;
	wire n579, n577, n580, n583, n973, n993, n1186, n584, n582, n1006, n585;
	wire n590, n588, n591, n594, n596, n601, n605, n611, n789, n1259, n612;
	wire n610, n689, n614, n1256, n615, n613, n1026, n617, n616, n619, n618;
	wire n623, n621, n626, n624, n628, n627, n630, n632, n633, n634, n638;
	wire n641, n644, n643, n642, n646, n645, n1004, n647, n1179, n651, n650;
	wire n653, n654, n652, n657, n655, n660, n1180, n1181, n1029, n661, n659;
	wire n658, n849, n665, n891, n668, n1024, n667, n672, n671, n1175, n676;
	wire n674, n677, n680, n682, n679, n683, n686, n691, n695, n696, n694;
	wire n1174, n698, n1021, n699, n697, n700, n1260, n703, n702, n705, n1022;
	wire n710, n709, n712, n714, n713, n718, n715, n720, n721, n719, n723;
	wire n722, n725, n727, n728, n726, n729, n1170, n731, n733, n739, n737;
	wire n741, n740, n743, n744, n975, n747, n1008, n745, n749, n748, n1182;
	wire n750, n754, n907, n755, n1198, n756, n1164, n1199, n1201, n757, n758;
	wire n759, n1202, n1172, n1203, n760, n1204, n1205, n1206, n1207, n1208, n1210;
	wire n761, n762, n764, n765, n767, n766, n951, n768, n771, n773, n777;
	wire n778, n776, n1242, n1241, n782, n781, n779, n1261, n784, n785, n783;
	wire n787, n790, n792, n791, n794, n793, n795, n797, n798, n796, n801;
	wire n799, n1040, n802, n806, n809, n810, n813, n812, n811, n824, n814;
	wire n818, n1272, n821, n828, n826, n823, n829, n1017, n1028, n827, n830;
	wire n831, n834, n837, n840, n843, n1043, n845, n847, n848, n851, n850;
	wire n1231, n868, n853, n1228, n854, n852, n855, n856, n857, n1276, n859;
	wire n1229, n861, n866, n1044, n864, n867, n870, n872, n871, n875, n873;
	wire n1038, n876, n882, n881, n883, n886, n1036, n888, n889, n887, n890;
	wire n892, n893, n895, n894, n897, n896, n898, n899, n901, n1279, n904;
	wire n906, n909, n908, n911, n910, n912, n1281, n916, n1216, n914, n931;
	wire n1257, n915, n913, n917, n919, n918, n920, n922, n921, n1039, n926;
	wire n924, n927, n929, n1280, n1223, n1224, n1227, n979, n998, n1002, n1018;
	wire n1019, n1041, n1042, n1050, n1056, n1060, n1068, n1070, n1072, n1071, n1073;
	wire n1074, n1076, n1079, n1082, n1083, n1084, n1085, n1087, n1092, n1094, n1100;
	wire n1099, n1101, n1107, n1109, n1112, n1127, n1120, n1122, n1124, n1128, n1130;
	wire n1131, n1134, n1133, n1135, n1136, n1140, n1226, n1264, n1147, n1155, n1171;
	wire n1173, n1183, n1189, n1191, n1195, n1197, n1200, n1268, n1209, n1214, n1222;
	wire n1220, n1225, n1230, n1232, n1237, n1236, n1238, n1239, n1244, n1243, n1245;
	wire n1247, n1246, n1273, n1251;



	assign o_0_ = (((!n1) & (!n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (!n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (!n3) & (n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (!n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (!n2) & (n3) & (n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (!n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (!n3) & (n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (!n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((!n1) & (n2) & (n3) & (n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((!n1) & (n2) & (n3) & (n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (!n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (!n3) & (n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (!n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (!n2) & (n3) & (n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (!n2) & (n3) & (n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (!n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (!n3) & (n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (!n3) & (n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (!n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (!n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (!n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (n3) & (!n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (!n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (!n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (n3) & (!n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (!n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (n3) & (!n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (!n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (n3) & (!n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (!n5) & (n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (n5) & (!n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (n3) & (n5) & (!n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (n5) & (!n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (n3) & (n5) & (!n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (n5) & (!n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (n3) & (n5) & (!n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (n5) & (!n8) & (n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (n3) & (n5) & (n8) & (!n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (n5) & (n8) & (!n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (n3) & (n5) & (n8) & (!n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (n5) & (n8) & (!n1248) & (n1249) & (n1250)) + ((n1) & (n2) & (n3) & (n5) & (n8) & (n1248) & (!n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (n5) & (n8) & (n1248) & (!n1249) & (n1250)) + ((n1) & (n2) & (n3) & (n5) & (n8) & (n1248) & (n1249) & (!n1250)) + ((n1) & (n2) & (n3) & (n5) & (n8) & (n1248) & (n1249) & (n1250)));
	assign o_1_ = (((!n753)));
	assign o_2_ = (((!n433)));
	assign n1 = (((n245) & (!n479) & (n880) & (!n1025)));
	assign n2 = (((i_35_) & (n670) & (n669) & (!n874)));
	assign n3 = (((!i_13_) & (!i_14_) & (!n885) & (!n1035)) + ((!i_13_) & (i_14_) & (!n885) & (!n1035)) + ((i_13_) & (!i_14_) & (!n885) & (!n1035)));
	assign n5 = (((!n216) & (!n608) & (!n662) & (!n1215)) + ((!n216) & (!n608) & (!n662) & (n1215)) + ((!n216) & (n608) & (!n662) & (!n1215)) + ((n216) & (!n608) & (!n662) & (!n1215)) + ((n216) & (n608) & (!n662) & (!n1215)));
	assign n8 = (((!n217) & (!n939) & (!n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (!n944) & (n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (!n942) & (n944) & (n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (!n944) & (n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (!n939) & (n942) & (n944) & (n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (!n944) & (n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (!n942) & (n944) & (n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (!n944) & (n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((!n217) & (n939) & (n942) & (n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((!n217) & (n939) & (n942) & (n944) & (n947) & (n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (!n944) & (n947) & (n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (!n942) & (n944) & (n947) & (n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (!n944) & (n947) & (n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (!n939) & (n942) & (n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (!n939) & (n942) & (n944) & (n947) & (n950) & (n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (!n944) & (n947) & (n950) & (n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (!n942) & (n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (!n942) & (n944) & (n947) & (n950) & (n1033) & (n1253)) + ((n217) & (n939) & (n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (!n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (n942) & (!n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (!n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (n939) & (n942) & (!n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (!n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (n942) & (!n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (!n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((n217) & (n939) & (n942) & (!n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (!n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (n942) & (!n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (!n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (n939) & (n942) & (!n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (!n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (n942) & (!n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (!n944) & (n947) & (n950) & (n1033) & (n1253)) + ((n217) & (n939) & (n942) & (n944) & (!n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (n944) & (!n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (n942) & (n944) & (!n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (n944) & (!n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (n939) & (n942) & (n944) & (!n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (n944) & (!n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (n942) & (n944) & (!n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (n944) & (!n947) & (n950) & (n1033) & (n1253)) + ((n217) & (n939) & (n942) & (n944) & (n947) & (!n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (n944) & (n947) & (!n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (n942) & (n944) & (n947) & (!n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (n944) & (n947) & (!n950) & (n1033) & (n1253)) + ((n217) & (n939) & (n942) & (n944) & (n947) & (n950) & (!n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (n944) & (n947) & (n950) & (!n1033) & (n1253)) + ((n217) & (n939) & (n942) & (n944) & (n947) & (n950) & (n1033) & (!n1253)) + ((n217) & (n939) & (n942) & (n944) & (n947) & (n950) & (n1033) & (n1253)));
	assign n10 = (((!i_27_) & (!n163)));
	assign n11 = (((!i_30_) & (n350)));
	assign n9 = (((i_36_) & (!n10) & (!n11) & (!n1213)) + ((i_36_) & (!n10) & (n11) & (!n1213)) + ((i_36_) & (n10) & (!n11) & (!n1213)) + ((i_36_) & (n10) & (n11) & (!n1213)) + ((i_36_) & (n10) & (n11) & (n1213)));
	assign n15 = (((!i_12_) & (!i_13_)));
	assign n13 = (((!i_7_) & (!n15) & (!n1030)) + ((!i_7_) & (n15) & (!n1030)) + ((!i_7_) & (n15) & (n1030)));
	assign n19 = (((!i_11_) & (!i_19_)));
	assign n17 = (((!i_24_) & (!n19) & (!n60) & (!n59)) + ((!i_24_) & (!n19) & (!n60) & (n59)) + ((!i_24_) & (n19) & (!n60) & (!n59)) + ((!i_24_) & (n19) & (!n60) & (n59)) + ((!i_24_) & (n19) & (n60) & (!n59)));
	assign n24 = (((!i_13_) & (i_18_) & (i_19_)));
	assign n23 = (((!i_13_) & (i_18_)));
	assign n22 = (((!i_11_) & (!i_22_) & (n24) & (!n23)) + ((!i_11_) & (!i_22_) & (n24) & (n23)) + ((i_11_) & (!i_22_) & (!n24) & (n23)) + ((i_11_) & (!i_22_) & (n24) & (!n23)) + ((i_11_) & (!i_22_) & (n24) & (n23)));
	assign n26 = (((!i_24_) & (!n19) & (!n67) & (!n66)) + ((!i_24_) & (!n19) & (!n67) & (n66)) + ((!i_24_) & (n19) & (!n67) & (!n66)) + ((!i_24_) & (n19) & (!n67) & (n66)) + ((!i_24_) & (n19) & (n67) & (!n66)));
	assign n30 = (((i_17_) & (i_12_)));
	assign n31 = (((i_14_) & (i_13_)));
	assign n29 = (((i_22_) & (!n30) & (n31)) + ((i_22_) & (n30) & (!n31)) + ((i_22_) & (n30) & (n31)));
	assign n33 = (((!i_10_) & (!i_24_)));
	assign n32 = (((!i_13_) & (!i_24_) & (n33) & (!n70)) + ((!i_13_) & (i_24_) & (n33) & (!n70)) + ((i_13_) & (!i_24_) & (!n33) & (!n70)) + ((i_13_) & (!i_24_) & (n33) & (!n70)) + ((i_13_) & (i_24_) & (n33) & (!n70)));
	assign n35 = (((!i_24_) & (!n30) & (n31)) + ((!i_24_) & (n30) & (!n31)) + ((!i_24_) & (n30) & (n31)));
	assign n38 = (((!i_1_) & (!n966) & (n769)) + ((!i_1_) & (n966) & (!n769)) + ((!i_1_) & (n966) & (n769)) + ((i_1_) & (!n966) & (!n769)) + ((i_1_) & (!n966) & (n769)) + ((i_1_) & (n966) & (!n769)) + ((i_1_) & (n966) & (n769)));
	assign n39 = (((!i_18_) & (!n256)) + ((!i_18_) & (n256)) + ((i_18_) & (!n256)));
	assign n40 = (((!i_6_) & (n97)) + ((i_6_) & (!n97)) + ((i_6_) & (n97)));
	assign n36 = (((!n38) & (!n39) & (n40) & (!n256)) + ((!n38) & (n39) & (!n40) & (!n256)) + ((!n38) & (n39) & (n40) & (!n256)) + ((n38) & (!n39) & (n40) & (!n256)) + ((n38) & (!n39) & (n40) & (n256)) + ((n38) & (n39) & (!n40) & (!n256)) + ((n38) & (n39) & (!n40) & (n256)) + ((n38) & (n39) & (n40) & (!n256)) + ((n38) & (n39) & (n40) & (n256)));
	assign n44 = (((i_11_) & (!i_13_)));
	assign n41 = (((!i_18_) & (n44) & (!n147) & (!n1000)) + ((!i_18_) & (n44) & (n147) & (!n1000)) + ((i_18_) & (n44) & (!n147) & (!n1000)) + ((i_18_) & (n44) & (!n147) & (n1000)) + ((i_18_) & (n44) & (n147) & (!n1000)));
	assign n48 = (((i_9_) & (n44)));
	assign n45 = (((!i_18_) & (!n38) & (!n40) & (n48)) + ((!i_18_) & (!n38) & (n40) & (n48)) + ((i_18_) & (!n38) & (!n40) & (n48)) + ((i_18_) & (!n38) & (n40) & (n48)) + ((i_18_) & (n38) & (!n40) & (n48)));
	assign n52 = (((!n324) & (!n394) & (!n800)) + ((!n324) & (!n394) & (n800)) + ((!n324) & (n394) & (!n800)) + ((!n324) & (n394) & (n800)) + ((n324) & (!n394) & (!n800)) + ((n324) & (!n394) & (n800)) + ((n324) & (n394) & (!n800)));
	assign n50 = (((!n394) & (!n968)) + ((!n394) & (n968)) + ((n394) & (n968)));
	assign n49 = (((n52) & (!n50) & (!n121)) + ((n52) & (n50) & (!n121)) + ((n52) & (n50) & (n121)));
	assign n56 = (((!n90) & (!n135) & (!n324)) + ((!n90) & (n135) & (!n324)) + ((!n90) & (n135) & (n324)) + ((n90) & (!n135) & (!n324)) + ((n90) & (!n135) & (n324)) + ((n90) & (n135) & (!n324)) + ((n90) & (n135) & (n324)));
	assign n53 = (((n56) & (!n121) & (!n290) & (!n402)) + ((n56) & (!n121) & (!n290) & (n402)) + ((n56) & (!n121) & (n290) & (!n402)) + ((n56) & (!n121) & (n290) & (n402)) + ((n56) & (n121) & (!n290) & (!n402)) + ((n56) & (n121) & (!n290) & (n402)) + ((n56) & (n121) & (n290) & (!n402)));
	assign n60 = (((!i_9_) & (!i_18_) & (n990)) + ((!i_9_) & (i_18_) & (!n990)) + ((!i_9_) & (i_18_) & (n990)) + ((i_9_) & (!i_18_) & (!n990)) + ((i_9_) & (!i_18_) & (n990)) + ((i_9_) & (i_18_) & (!n990)) + ((i_9_) & (i_18_) & (n990)));
	assign n59 = (((!n371) & (n84)) + ((n371) & (!n84)) + ((n371) & (n84)));
	assign n57 = (((!n19) & (n60) & (!n59)) + ((!n19) & (n60) & (n59)) + ((n19) & (n60) & (n59)));
	assign n64 = (((!i_6_) & (!n964) & (n97)) + ((!i_6_) & (n964) & (!n97)) + ((!i_6_) & (n964) & (n97)) + ((i_6_) & (!n964) & (!n97)) + ((i_6_) & (!n964) & (n97)) + ((i_6_) & (n964) & (!n97)) + ((i_6_) & (n964) & (n97)));
	assign n63 = (((!n374) & (n965)) + ((n374) & (!n965)) + ((n374) & (n965)));
	assign n61 = (((!i_9_) & (n64) & (!n63)) + ((!i_9_) & (n64) & (n63)) + ((i_9_) & (n64) & (n63)));
	assign n67 = (((!i_18_) & (n985)) + ((i_18_) & (!n985)) + ((i_18_) & (n985)));
	assign n66 = (((!n371) & (n81)) + ((n371) & (!n81)) + ((n371) & (n81)));
	assign n65 = (((!n19) & (n67) & (!n66)) + ((!n19) & (n67) & (n66)) + ((n19) & (n67) & (n66)));
	assign n69 = (((i_10_) & (!i_13_)));
	assign n70 = (((!i_9_) & (n986)) + ((i_9_) & (!n986)) + ((i_9_) & (n986)));
	assign n68 = (((!n69) & (n70) & (!i_32_) & (n65)) + ((!n69) & (n70) & (i_32_) & (!n65)) + ((!n69) & (n70) & (i_32_) & (n65)) + ((n69) & (!n70) & (!i_32_) & (n65)) + ((n69) & (!n70) & (i_32_) & (!n65)) + ((n69) & (!n70) & (i_32_) & (n65)) + ((n69) & (n70) & (!i_32_) & (n65)) + ((n69) & (n70) & (i_32_) & (!n65)) + ((n69) & (n70) & (i_32_) & (n65)));
	assign n72 = (((!i_9_) & (!n965) & (!n977)) + ((!i_9_) & (!n965) & (n977)) + ((!i_9_) & (n965) & (!n977)) + ((!i_9_) & (n965) & (n977)) + ((i_9_) & (!n965) & (n977)) + ((i_9_) & (n965) & (!n977)) + ((i_9_) & (n965) & (n977)));
	assign n73 = (((!i_11_) & (!i_12_)) + ((!i_11_) & (i_12_)) + ((i_11_) & (i_12_)));
	assign n74 = (((!i_11_) & (!n964)) + ((!i_11_) & (n964)) + ((i_11_) & (n964)));
	assign n71 = (((!n72) & (n73) & (!n38) & (n74)) + ((!n72) & (n73) & (n38) & (!n74)) + ((!n72) & (n73) & (n38) & (n74)) + ((n72) & (!n73) & (!n38) & (n74)) + ((n72) & (!n73) & (n38) & (!n74)) + ((n72) & (!n73) & (n38) & (n74)) + ((n72) & (n73) & (!n38) & (n74)) + ((n72) & (n73) & (n38) & (!n74)) + ((n72) & (n73) & (n38) & (n74)));
	assign n75 = (((!n44) & (!n48) & (!n64) & (!n63)) + ((!n44) & (!n48) & (!n64) & (n63)) + ((!n44) & (!n48) & (n64) & (!n63)) + ((!n44) & (!n48) & (n64) & (n63)) + ((!n44) & (n48) & (!n64) & (n63)) + ((!n44) & (n48) & (n64) & (n63)) + ((n44) & (!n48) & (n64) & (!n63)) + ((n44) & (!n48) & (n64) & (n63)) + ((n44) & (n48) & (n64) & (n63)));
	assign n78 = (((!i_13_) & (!i_18_) & (n71) & (!n75)) + ((!i_13_) & (!i_18_) & (n71) & (n75)) + ((!i_13_) & (i_18_) & (n71) & (n75)) + ((i_13_) & (!i_18_) & (!n71) & (!n75)) + ((i_13_) & (!i_18_) & (!n71) & (n75)) + ((i_13_) & (!i_18_) & (n71) & (!n75)) + ((i_13_) & (!i_18_) & (n71) & (n75)) + ((i_13_) & (i_18_) & (!n71) & (n75)) + ((i_13_) & (i_18_) & (n71) & (n75)));
	assign n81 = (((!i_7_) & (n989)) + ((i_7_) & (!n989)) + ((i_7_) & (n989)));
	assign n82 = (((!i_32_) & (!i_38_)) + ((i_32_) & (!i_38_)) + ((i_32_) & (i_38_)));
	assign n84 = (((!i_8_) & (n989)) + ((i_8_) & (!n989)) + ((i_8_) & (n989)));
	assign n80 = (((!n81) & (n82) & (!n84) & (!n299)) + ((!n81) & (n82) & (n84) & (!n299)) + ((!n81) & (n82) & (n84) & (n299)) + ((n81) & (!n82) & (!n84) & (!n299)) + ((n81) & (!n82) & (n84) & (!n299)) + ((n81) & (!n82) & (n84) & (n299)) + ((n81) & (n82) & (!n84) & (!n299)) + ((n81) & (n82) & (n84) & (!n299)) + ((n81) & (n82) & (n84) & (n299)));
	assign n87 = (((!n81) & (!n91) & (!n322)) + ((!n81) & (n91) & (!n322)) + ((!n81) & (n91) & (n322)) + ((n81) & (!n91) & (!n322)) + ((n81) & (!n91) & (n322)) + ((n81) & (n91) & (!n322)) + ((n81) & (n91) & (n322)));
	assign n88 = (((!n84) & (!n100) & (!n402)) + ((!n84) & (n100) & (!n402)) + ((!n84) & (n100) & (n402)) + ((n84) & (!n100) & (!n402)) + ((n84) & (!n100) & (n402)) + ((n84) & (n100) & (!n402)) + ((n84) & (n100) & (n402)));
	assign n86 = (((!i_25_) & (n963)) + ((i_25_) & (!n963)) + ((i_25_) & (n963)));
	assign n85 = (((n87) & (n88) & (!n80) & (n86)) + ((n87) & (n88) & (n80) & (!n86)) + ((n87) & (n88) & (n80) & (n86)));
	assign n90 = (((!i_32_) & (!n394)) + ((i_32_) & (!n394)) + ((i_32_) & (n394)));
	assign n91 = (((!i_32_) & (n963)) + ((i_32_) & (!n963)) + ((i_32_) & (n963)));
	assign n89 = (((!n86) & (n90) & (!n91) & (!n402)) + ((!n86) & (n90) & (n91) & (!n402)) + ((!n86) & (n90) & (n91) & (n402)) + ((n86) & (!n90) & (!n91) & (!n402)) + ((n86) & (!n90) & (n91) & (!n402)) + ((n86) & (!n90) & (n91) & (n402)) + ((n86) & (n90) & (!n91) & (!n402)) + ((n86) & (n90) & (n91) & (!n402)) + ((n86) & (n90) & (n91) & (n402)));
	assign n93 = (((!n983) & (n528)) + ((n983) & (!n528)) + ((n983) & (n528)));
	assign n94 = (((!n371) & (n991)) + ((n371) & (!n991)) + ((n371) & (n991)));
	assign n92 = (((!i_18_) & (n93) & (!i_19_) & (n94)) + ((!i_18_) & (n93) & (i_19_) & (!n94)) + ((!i_18_) & (n93) & (i_19_) & (n94)) + ((i_18_) & (!n93) & (!i_19_) & (n94)) + ((i_18_) & (!n93) & (i_19_) & (!n94)) + ((i_18_) & (!n93) & (i_19_) & (n94)) + ((i_18_) & (n93) & (!i_19_) & (n94)) + ((i_18_) & (n93) & (i_19_) & (!n94)) + ((i_18_) & (n93) & (i_19_) & (n94)));
	assign n96 = (((!n374) & (n595)) + ((n374) & (!n595)) + ((n374) & (n595)));
	assign n97 = (((!i_12_) & (n371)) + ((i_12_) & (!n371)) + ((i_12_) & (n371)));
	assign n98 = (((!i_6_) & (!n229)) + ((i_6_) & (!n229)) + ((i_6_) & (n229)));
	assign n95 = (((!i_8_) & (n96) & (!n97) & (n98)) + ((!i_8_) & (n96) & (n97) & (!n98)) + ((!i_8_) & (n96) & (n97) & (n98)) + ((i_8_) & (!n96) & (!n97) & (n98)) + ((i_8_) & (!n96) & (n97) & (!n98)) + ((i_8_) & (!n96) & (n97) & (n98)) + ((i_8_) & (n96) & (!n97) & (n98)) + ((i_8_) & (n96) & (n97) & (!n98)) + ((i_8_) & (n96) & (n97) & (n98)));
	assign n100 = (((!i_31_) & (n963)) + ((i_31_) & (!n963)) + ((i_31_) & (n963)));
	assign n101 = (((!i_35_) & (n970)) + ((i_35_) & (!n970)) + ((i_35_) & (n970)));
	assign n99 = (((!n100) & (!n92) & (n101)) + ((!n100) & (n92) & (!n101)) + ((!n100) & (n92) & (n101)) + ((n100) & (!n92) & (!n101)) + ((n100) & (!n92) & (n101)) + ((n100) & (n92) & (!n101)) + ((n100) & (n92) & (n101)));
	assign n104 = (((!i_32_) & (!n92) & (!n299)) + ((!i_32_) & (n92) & (!n299)) + ((!i_32_) & (n92) & (n299)) + ((i_32_) & (!n92) & (!n299)) + ((i_32_) & (!n92) & (n299)) + ((i_32_) & (n92) & (!n299)) + ((i_32_) & (n92) & (n299)));
	assign n102 = (((!i_2_) & (n104) & (!n290) & (!n394)) + ((!i_2_) & (n104) & (!n290) & (n394)) + ((!i_2_) & (n104) & (n290) & (!n394)) + ((i_2_) & (n104) & (!n290) & (!n394)) + ((i_2_) & (n104) & (!n290) & (n394)) + ((i_2_) & (n104) & (n290) & (!n394)) + ((i_2_) & (n104) & (n290) & (n394)));
	assign n107 = (((!n86) & (!n1258)) + ((!n86) & (n1258)) + ((n86) & (!n1258)));
	assign n105 = (((i_38_) & (!n95) & (!n99) & (!n107)) + ((i_38_) & (!n95) & (!n99) & (n107)) + ((i_38_) & (!n95) & (n99) & (n107)) + ((i_38_) & (n95) & (!n99) & (!n107)) + ((i_38_) & (n95) & (!n99) & (n107)));
	assign n112 = (((!n800) & (!n1001) & (n1117)) + ((!n800) & (n1001) & (n1117)) + ((n800) & (n1001) & (n1117)));
	assign n110 = (((!i_38_) & (!n57) & (!n68) & (!n299)) + ((!i_38_) & (!n57) & (n68) & (!n299)) + ((!i_38_) & (n57) & (!n68) & (!n299)) + ((!i_38_) & (n57) & (!n68) & (n299)) + ((!i_38_) & (n57) & (n68) & (!n299)) + ((!i_38_) & (n57) & (n68) & (n299)) + ((i_38_) & (!n57) & (n68) & (!n299)) + ((i_38_) & (n57) & (n68) & (!n299)) + ((i_38_) & (n57) & (n68) & (n299)));
	assign n111 = (((!i_10_) & (!n61) & (!n394) & (n1116)) + ((!i_10_) & (n61) & (!n394) & (n1116)) + ((!i_10_) & (n61) & (n394) & (n1116)) + ((i_10_) & (!n61) & (!n394) & (n1116)) + ((i_10_) & (!n61) & (n394) & (n1116)) + ((i_10_) & (n61) & (!n394) & (n1116)) + ((i_10_) & (n61) & (n394) & (n1116)));
	assign n109 = (((n112) & (!i_28_) & (n110) & (n111)) + ((n112) & (i_28_) & (!n110) & (!n111)) + ((n112) & (i_28_) & (!n110) & (n111)) + ((n112) & (i_28_) & (n110) & (!n111)) + ((n112) & (i_28_) & (n110) & (n111)));
	assign n113 = (((!i_24_) & (!n1118) & (!n1121) & (!n1123)) + ((!i_24_) & (!n1118) & (!n1121) & (n1123)) + ((!i_24_) & (!n1118) & (n1121) & (!n1123)) + ((!i_24_) & (!n1118) & (n1121) & (n1123)) + ((!i_24_) & (n1118) & (!n1121) & (!n1123)) + ((!i_24_) & (n1118) & (!n1121) & (n1123)) + ((!i_24_) & (n1118) & (n1121) & (!n1123)));
	assign n121 = (((!i_28_) & (!n163)));
	assign n117 = (((n121) & (!n1126) & (!n1129) & (!n1132)) + ((n121) & (!n1126) & (!n1129) & (n1132)) + ((n121) & (!n1126) & (n1129) & (!n1132)) + ((n121) & (!n1126) & (n1129) & (n1132)) + ((n121) & (n1126) & (!n1129) & (!n1132)) + ((n121) & (n1126) & (!n1129) & (n1132)) + ((n121) & (n1126) & (n1129) & (!n1132)));
	assign n125 = (((!i_30_) & (!n162) & (!n313)) + ((!i_30_) & (n162) & (!n313)) + ((!i_30_) & (n162) & (n313)) + ((i_30_) & (!n162) & (!n313)) + ((i_30_) & (!n162) & (n313)) + ((i_30_) & (n162) & (!n313)) + ((i_30_) & (n162) & (n313)));
	assign n126 = (((!n86) & (!n195) & (!n306) & (n994)) + ((!n86) & (n195) & (!n306) & (n994)) + ((!n86) & (n195) & (n306) & (n994)) + ((n86) & (!n195) & (!n306) & (!n994)) + ((n86) & (!n195) & (!n306) & (n994)) + ((n86) & (n195) & (!n306) & (!n994)) + ((n86) & (n195) & (!n306) & (n994)) + ((n86) & (n195) & (n306) & (!n994)) + ((n86) & (n195) & (n306) & (n994)));
	assign n124 = (((!i_38_) & (!n988)) + ((!i_38_) & (n988)) + ((i_38_) & (n988)));
	assign n122 = (((!n11) & (n125) & (n126) & (!n124)) + ((!n11) & (n125) & (n126) & (n124)) + ((n11) & (n125) & (n126) & (n124)));
	assign n129 = (((!i_28_) & (n179)) + ((i_28_) & (!n179)) + ((i_28_) & (n179)));
	assign n130 = (((!i_22_) & (!n288)) + ((i_22_) & (!n288)) + ((i_22_) & (n288)));
	assign n131 = (((!n138) & (!n394)) + ((n138) & (!n394)) + ((n138) & (n394)));
	assign n127 = (((!n129) & (!n130) & (n131) & (!n306)) + ((!n129) & (n130) & (!n131) & (!n306)) + ((!n129) & (n130) & (n131) & (!n306)) + ((n129) & (!n130) & (n131) & (!n306)) + ((n129) & (!n130) & (n131) & (n306)) + ((n129) & (n130) & (!n131) & (!n306)) + ((n129) & (n130) & (!n131) & (n306)) + ((n129) & (n130) & (n131) & (!n306)) + ((n129) & (n130) & (n131) & (n306)));
	assign n133 = (((!n130) & (n138)) + ((n130) & (!n138)) + ((n130) & (n138)));
	assign n134 = (((!n179) & (!n402)) + ((n179) & (!n402)) + ((n179) & (n402)));
	assign n135 = (((!i_31_) & (!i_30_) & (i_28_)) + ((!i_31_) & (i_30_) & (!i_28_)) + ((!i_31_) & (i_30_) & (i_28_)) + ((i_31_) & (!i_30_) & (!i_28_)) + ((i_31_) & (!i_30_) & (i_28_)) + ((i_31_) & (i_30_) & (!i_28_)) + ((i_31_) & (i_30_) & (i_28_)));
	assign n132 = (((!n133) & (!n134) & (n135) & (!n299)) + ((!n133) & (n134) & (!n135) & (!n299)) + ((!n133) & (n134) & (n135) & (!n299)) + ((n133) & (!n134) & (n135) & (!n299)) + ((n133) & (!n134) & (n135) & (n299)) + ((n133) & (n134) & (!n135) & (!n299)) + ((n133) & (n134) & (!n135) & (n299)) + ((n133) & (n134) & (n135) & (!n299)) + ((n133) & (n134) & (n135) & (n299)));
	assign n139 = (((!i_30_) & (!i_38_) & (!n86)) + ((!i_30_) & (!i_38_) & (n86)) + ((!i_30_) & (i_38_) & (n86)) + ((i_30_) & (!i_38_) & (!n86)) + ((i_30_) & (!i_38_) & (n86)) + ((i_30_) & (i_38_) & (!n86)) + ((i_30_) & (i_38_) & (n86)));
	assign n138 = (((!i_30_) & (n963)) + ((i_30_) & (!n963)) + ((i_30_) & (n963)));
	assign n136 = (((n139) & (!n138) & (!n322)) + ((n139) & (n138) & (!n322)) + ((n139) & (n138) & (n322)));
	assign n140 = (((!n33) & (!n64) & (!n63) & (!n311)) + ((!n33) & (!n64) & (n63) & (!n311)) + ((!n33) & (!n64) & (n63) & (n311)) + ((!n33) & (n64) & (!n63) & (!n311)) + ((!n33) & (n64) & (n63) & (!n311)) + ((!n33) & (n64) & (n63) & (n311)) + ((n33) & (n64) & (!n63) & (!n311)) + ((n33) & (n64) & (n63) & (!n311)) + ((n33) & (n64) & (n63) & (n311)));
	assign n144 = (((!i_18_) & (!n288)) + ((!i_18_) & (n288)) + ((i_18_) & (!n288)));
	assign n145 = (((!i_13_) & (!n288)) + ((i_13_) & (!n288)) + ((i_13_) & (n288)));
	assign n143 = (((!n75) & (n144) & (!n71) & (n145)) + ((!n75) & (n144) & (n71) & (!n145)) + ((!n75) & (n144) & (n71) & (n145)) + ((n75) & (!n144) & (!n71) & (n145)) + ((n75) & (!n144) & (n71) & (!n145)) + ((n75) & (!n144) & (n71) & (n145)) + ((n75) & (n144) & (!n71) & (n145)) + ((n75) & (n144) & (n71) & (!n145)) + ((n75) & (n144) & (n71) & (n145)));
	assign n147 = (((!n962) & (n374)) + ((n962) & (!n374)) + ((n962) & (n374)));
	assign n148 = (((!i_6_) & (!i_9_) & (!i_10_)) + ((!i_6_) & (!i_9_) & (i_10_)) + ((!i_6_) & (i_9_) & (i_10_)) + ((i_6_) & (!i_9_) & (!i_10_)) + ((i_6_) & (!i_9_) & (i_10_)) + ((i_6_) & (i_9_) & (!i_10_)) + ((i_6_) & (i_9_) & (i_10_)));
	assign n146 = (((!i_10_) & (n147) & (!n97) & (n148)) + ((!i_10_) & (n147) & (n97) & (!n148)) + ((!i_10_) & (n147) & (n97) & (n148)) + ((i_10_) & (!n147) & (!n97) & (n148)) + ((i_10_) & (!n147) & (n97) & (!n148)) + ((i_10_) & (!n147) & (n97) & (n148)) + ((i_10_) & (n147) & (!n97) & (n148)) + ((i_10_) & (n147) & (n97) & (!n148)) + ((i_10_) & (n147) & (n97) & (n148)));
	assign n150 = (((!i_8_) & (!i_30_) & (!n299)) + ((!i_8_) & (i_30_) & (!n299)) + ((!i_8_) & (i_30_) & (n299)) + ((i_8_) & (!i_30_) & (!n299)) + ((i_8_) & (!i_30_) & (n299)) + ((i_8_) & (i_30_) & (!n299)) + ((i_8_) & (i_30_) & (n299)));
	assign n151 = (((n104) & (!n69) & (!n80) & (n371)) + ((n104) & (!n69) & (n80) & (!n371)) + ((n104) & (!n69) & (n80) & (n371)) + ((n104) & (n69) & (!n80) & (!n371)) + ((n104) & (n69) & (!n80) & (n371)) + ((n104) & (n69) & (n80) & (!n371)) + ((n104) & (n69) & (n80) & (n371)));
	assign n149 = (((n150) & (n151) & (!n146) & (n90)) + ((n150) & (n151) & (n146) & (!n90)) + ((n150) & (n151) & (n146) & (n90)));
	assign n152 = (((!i_32_) & (!n26) & (!n32)) + ((i_32_) & (!n26) & (!n32)) + ((i_32_) & (n26) & (!n32)));
	assign n155 = (((!i_30_) & (n152) & (!n414)) + ((i_30_) & (n152) & (!n414)) + ((i_30_) & (n152) & (n414)));
	assign n159 = (((!n17) & (!n155) & (!n322) & (!n326)) + ((!n17) & (!n155) & (!n322) & (n326)) + ((!n17) & (n155) & (!n322) & (!n326)) + ((!n17) & (n155) & (!n322) & (n326)) + ((!n17) & (n155) & (n322) & (!n326)) + ((!n17) & (n155) & (n322) & (n326)) + ((n17) & (!n155) & (!n322) & (n326)) + ((n17) & (n155) & (!n322) & (n326)) + ((n17) & (n155) & (n322) & (n326)));
	assign n160 = (((!n50) & (!n311) & (n1115)) + ((n50) & (!n311) & (n1115)) + ((n50) & (n311) & (n1115)));
	assign n157 = (((!n149) & (n159) & (n160) & (!n288)) + ((n149) & (n159) & (n160) & (!n288)) + ((n149) & (n159) & (n160) & (n288)));
	assign n162 = (((!i_34_) & (!n394)) + ((!i_34_) & (n394)) + ((i_34_) & (!n394)));
	assign n163 = (((!i_24_) & (i_26_)) + ((i_24_) & (!i_26_)) + ((i_24_) & (i_26_)));
	assign n161 = (((!n162) & (!n163) & (!n288) & (!n402)) + ((!n162) & (n163) & (!n288) & (!n402)) + ((!n162) & (n163) & (!n288) & (n402)) + ((n162) & (!n163) & (!n288) & (!n402)) + ((n162) & (!n163) & (n288) & (!n402)) + ((n162) & (n163) & (!n288) & (!n402)) + ((n162) & (n163) & (!n288) & (n402)) + ((n162) & (n163) & (n288) & (!n402)) + ((n162) & (n163) & (n288) & (n402)));
	assign n167 = (((!n81) & (!n163) & (!n322) & (!n367)) + ((!n81) & (!n163) & (!n322) & (n367)) + ((!n81) & (!n163) & (n322) & (!n367)) + ((!n81) & (n163) & (!n322) & (!n367)) + ((!n81) & (n163) & (!n322) & (n367)) + ((!n81) & (n163) & (n322) & (!n367)) + ((!n81) & (n163) & (n322) & (n367)) + ((n81) & (!n163) & (!n322) & (!n367)) + ((n81) & (!n163) & (!n322) & (n367)) + ((n81) & (!n163) & (n322) & (!n367)) + ((n81) & (!n163) & (n322) & (n367)) + ((n81) & (n163) & (!n322) & (!n367)) + ((n81) & (n163) & (!n322) & (n367)) + ((n81) & (n163) & (n322) & (!n367)) + ((n81) & (n163) & (n322) & (n367)));
	assign n165 = (((!n161) & (n170)) + ((n161) & (!n170)) + ((n161) & (n170)));
	assign n166 = (((!i_31_) & (!i_33_) & (!n162) & (!n308)) + ((!i_31_) & (!i_33_) & (n162) & (!n308)) + ((!i_31_) & (!i_33_) & (n162) & (n308)) + ((!i_31_) & (i_33_) & (!n162) & (!n308)) + ((!i_31_) & (i_33_) & (!n162) & (n308)) + ((!i_31_) & (i_33_) & (n162) & (!n308)) + ((!i_31_) & (i_33_) & (n162) & (n308)) + ((i_31_) & (!i_33_) & (!n162) & (!n308)) + ((i_31_) & (!i_33_) & (!n162) & (n308)) + ((i_31_) & (!i_33_) & (n162) & (!n308)) + ((i_31_) & (!i_33_) & (n162) & (n308)) + ((i_31_) & (i_33_) & (!n162) & (!n308)) + ((i_31_) & (i_33_) & (!n162) & (n308)) + ((i_31_) & (i_33_) & (n162) & (!n308)) + ((i_31_) & (i_33_) & (n162) & (n308)));
	assign n164 = (((n167) & (!n84) & (n165) & (n166)) + ((n167) & (n84) & (!n165) & (!n166)) + ((n167) & (n84) & (!n165) & (n166)) + ((n167) & (n84) & (n165) & (!n166)) + ((n167) & (n84) & (n165) & (n166)));
	assign n170 = (((!i_31_) & (!n350)) + ((i_31_) & (!n350)) + ((i_31_) & (n350)));
	assign n168 = (((!n100) & (n130) & (!n170) & (!n324)) + ((!n100) & (n130) & (n170) & (!n324)) + ((!n100) & (n130) & (n170) & (n324)) + ((n100) & (!n130) & (!n170) & (!n324)) + ((n100) & (!n130) & (n170) & (!n324)) + ((n100) & (!n130) & (n170) & (n324)) + ((n100) & (n130) & (!n170) & (!n324)) + ((n100) & (n130) & (n170) & (!n324)) + ((n100) & (n130) & (n170) & (n324)));
	assign n171 = (((!n121) & (!n162) & (!n304) & (!n402)) + ((!n121) & (!n162) & (!n304) & (n402)) + ((!n121) & (n162) & (!n304) & (!n402)) + ((!n121) & (n162) & (!n304) & (n402)) + ((!n121) & (n162) & (n304) & (!n402)) + ((!n121) & (n162) & (n304) & (n402)) + ((n121) & (!n162) & (!n304) & (!n402)) + ((n121) & (n162) & (!n304) & (!n402)) + ((n121) & (n162) & (n304) & (!n402)));
	assign n175 = (((!n162) & (!n308) & (!n972)) + ((!n162) & (!n308) & (n972)) + ((!n162) & (n308) & (n972)) + ((n162) & (!n308) & (!n972)) + ((n162) & (!n308) & (n972)) + ((n162) & (n308) & (!n972)) + ((n162) & (n308) & (n972)));
	assign n176 = (((!n168) & (n90) & (!i_31_) & (n206)) + ((!n168) & (n90) & (i_31_) & (!n206)) + ((!n168) & (n90) & (i_31_) & (n206)) + ((n168) & (!n90) & (!i_31_) & (n206)) + ((n168) & (!n90) & (i_31_) & (!n206)) + ((n168) & (!n90) & (i_31_) & (n206)) + ((n168) & (n90) & (!i_31_) & (n206)) + ((n168) & (n90) & (i_31_) & (!n206)) + ((n168) & (n90) & (i_31_) & (n206)));
	assign n174 = (((!i_29_) & (n685)) + ((i_29_) & (!n685)) + ((i_29_) & (n685)));
	assign n173 = (((n175) & (n176) & (!n171) & (n174)) + ((n175) & (n176) & (n171) & (!n174)) + ((n175) & (n176) & (n171) & (n174)));
	assign n180 = (((!i_32_) & (!i_38_) & (!n130) & (!n138)) + ((!i_32_) & (!i_38_) & (!n130) & (n138)) + ((!i_32_) & (!i_38_) & (n130) & (!n138)) + ((!i_32_) & (!i_38_) & (n130) & (n138)) + ((!i_32_) & (i_38_) & (!n130) & (n138)) + ((!i_32_) & (i_38_) & (n130) & (!n138)) + ((!i_32_) & (i_38_) & (n130) & (n138)) + ((i_32_) & (!i_38_) & (!n130) & (!n138)) + ((i_32_) & (!i_38_) & (!n130) & (n138)) + ((i_32_) & (!i_38_) & (n130) & (!n138)) + ((i_32_) & (!i_38_) & (n130) & (n138)) + ((i_32_) & (i_38_) & (!n130) & (!n138)) + ((i_32_) & (i_38_) & (!n130) & (n138)) + ((i_32_) & (i_38_) & (n130) & (!n138)) + ((i_32_) & (i_38_) & (n130) & (n138)));
	assign n179 = (((!i_22_) & (n163)) + ((i_22_) & (!n163)) + ((i_22_) & (n163)));
	assign n177 = (((n180) & (!n179) & (!n322) & (!n800)) + ((n180) & (!n179) & (!n322) & (n800)) + ((n180) & (!n179) & (n322) & (!n800)) + ((n180) & (n179) & (!n322) & (!n800)) + ((n180) & (n179) & (!n322) & (n800)) + ((n180) & (n179) & (n322) & (!n800)) + ((n180) & (n179) & (n322) & (n800)));
	assign n183 = (((!n177) & (n987)) + ((n177) & (!n987)) + ((n177) & (n987)));
	assign n184 = (((!i_3_) & (!i_8_) & (!i_10_) & (!n132)) + ((!i_3_) & (!i_8_) & (!i_10_) & (n132)) + ((!i_3_) & (!i_8_) & (i_10_) & (n132)) + ((!i_3_) & (i_8_) & (!i_10_) & (!n132)) + ((!i_3_) & (i_8_) & (!i_10_) & (n132)) + ((!i_3_) & (i_8_) & (i_10_) & (!n132)) + ((!i_3_) & (i_8_) & (i_10_) & (n132)) + ((i_3_) & (!i_8_) & (!i_10_) & (!n132)) + ((i_3_) & (!i_8_) & (!i_10_) & (n132)) + ((i_3_) & (!i_8_) & (i_10_) & (!n132)) + ((i_3_) & (!i_8_) & (i_10_) & (n132)) + ((i_3_) & (i_8_) & (!i_10_) & (!n132)) + ((i_3_) & (i_8_) & (!i_10_) & (n132)) + ((i_3_) & (i_8_) & (i_10_) & (!n132)) + ((i_3_) & (i_8_) & (i_10_) & (n132)));
	assign n182 = (((!i_3_) & (n964)) + ((i_3_) & (!n964)) + ((i_3_) & (n964)));
	assign n181 = (((n183) & (n184) & (!n127) & (n182)) + ((n183) & (n184) & (n127) & (!n182)) + ((n183) & (n184) & (n127) & (n182)));
	assign n185 = (((!i_28_) & (!i_29_) & (!n121) & (n179)) + ((!i_28_) & (i_29_) & (!n121) & (n179)) + ((!i_28_) & (i_29_) & (n121) & (n179)) + ((i_28_) & (!i_29_) & (!n121) & (!n179)) + ((i_28_) & (!i_29_) & (!n121) & (n179)) + ((i_28_) & (i_29_) & (!n121) & (!n179)) + ((i_28_) & (i_29_) & (!n121) & (n179)) + ((i_28_) & (i_29_) & (n121) & (!n179)) + ((i_28_) & (i_29_) & (n121) & (n179)));
	assign n188 = (((!i_2_) & (n964)) + ((i_2_) & (!n964)) + ((i_2_) & (n964)));
	assign n189 = (((!i_12_) & (!i_22_) & (!i_24_)) + ((!i_12_) & (!i_22_) & (i_24_)) + ((!i_12_) & (i_22_) & (!i_24_)) + ((!i_12_) & (i_22_) & (i_24_)) + ((i_12_) & (!i_22_) & (i_24_)) + ((i_12_) & (i_22_) & (!i_24_)) + ((i_12_) & (i_22_) & (i_24_)));
	assign n190 = (((!i_10_) & (n964)) + ((i_10_) & (!n964)) + ((i_10_) & (n964)));
	assign n186 = (((!n188) & (!n189) & (n190) & (!n429)) + ((!n188) & (n189) & (!n190) & (!n429)) + ((!n188) & (n189) & (n190) & (!n429)) + ((n188) & (!n189) & (n190) & (!n429)) + ((n188) & (!n189) & (n190) & (n429)) + ((n188) & (n189) & (!n190) & (!n429)) + ((n188) & (n189) & (!n190) & (n429)) + ((n188) & (n189) & (n190) & (!n429)) + ((n188) & (n189) & (n190) & (n429)));
	assign n193 = (((!i_26_) & (!i_38_) & (!n11) & (!n101)) + ((!i_26_) & (!i_38_) & (!n11) & (n101)) + ((!i_26_) & (!i_38_) & (n11) & (!n101)) + ((!i_26_) & (!i_38_) & (n11) & (n101)) + ((!i_26_) & (i_38_) & (!n11) & (!n101)) + ((!i_26_) & (i_38_) & (!n11) & (n101)) + ((!i_26_) & (i_38_) & (n11) & (n101)) + ((i_26_) & (!i_38_) & (!n11) & (!n101)) + ((i_26_) & (!i_38_) & (!n11) & (n101)) + ((i_26_) & (!i_38_) & (n11) & (!n101)) + ((i_26_) & (!i_38_) & (n11) & (n101)) + ((i_26_) & (i_38_) & (!n11) & (!n101)) + ((i_26_) & (i_38_) & (!n11) & (n101)) + ((i_26_) & (i_38_) & (n11) & (!n101)) + ((i_26_) & (i_38_) & (n11) & (n101)));
	assign n192 = (((!i_29_) & (!n234)) + ((i_29_) & (!n234)) + ((i_29_) & (n234)));
	assign n191 = (((n193) & (!i_28_) & (!n192) & (n124)) + ((n193) & (!i_28_) & (n192) & (!n124)) + ((n193) & (!i_28_) & (n192) & (n124)) + ((n193) & (i_28_) & (!n192) & (!n124)) + ((n193) & (i_28_) & (!n192) & (n124)) + ((n193) & (i_28_) & (n192) & (!n124)) + ((n193) & (i_28_) & (n192) & (n124)));
	assign n197 = (((!i_38_) & (!n11) & (!n832)) + ((!i_38_) & (!n11) & (n832)) + ((!i_38_) & (n11) & (!n832)) + ((!i_38_) & (n11) & (n832)) + ((i_38_) & (!n11) & (!n832)) + ((i_38_) & (!n11) & (n832)) + ((i_38_) & (n11) & (!n832)));
	assign n195 = (((!i_26_) & (!n350)) + ((i_26_) & (!n350)) + ((i_26_) & (n350)));
	assign n196 = (((!i_30_) & (n90)) + ((i_30_) & (!n90)) + ((i_30_) & (n90)));
	assign n194 = (((n197) & (!n195) & (n196)) + ((n197) & (n195) & (!n196)) + ((n197) & (n195) & (n196)));
	assign n199 = (((!i_19_) & (!i_24_)) + ((!i_19_) & (i_24_)) + ((i_19_) & (i_24_)));
	assign n200 = (((!i_19_) & (!n288)) + ((!i_19_) & (n288)) + ((i_19_) & (!n288)));
	assign n198 = (((!n191) & (n199) & (!n194) & (n200)) + ((!n191) & (n199) & (n194) & (!n200)) + ((!n191) & (n199) & (n194) & (n200)) + ((n191) & (!n199) & (!n194) & (n200)) + ((n191) & (!n199) & (n194) & (!n200)) + ((n191) & (!n199) & (n194) & (n200)) + ((n191) & (n199) & (!n194) & (n200)) + ((n191) & (n199) & (n194) & (!n200)) + ((n191) & (n199) & (n194) & (n200)));
	assign n203 = (((!n91) & (n130) & (!n304) & (!n648)) + ((!n91) & (n130) & (!n304) & (n648)) + ((!n91) & (n130) & (n304) & (n648)) + ((n91) & (!n130) & (!n304) & (!n648)) + ((n91) & (!n130) & (!n304) & (n648)) + ((n91) & (!n130) & (n304) & (n648)) + ((n91) & (n130) & (!n304) & (!n648)) + ((n91) & (n130) & (!n304) & (n648)) + ((n91) & (n130) & (n304) & (n648)));
	assign n204 = (((!n121) & (!n241) & (!n308) & (!n376)) + ((!n121) & (!n241) & (!n308) & (n376)) + ((!n121) & (!n241) & (n308) & (n376)) + ((!n121) & (n241) & (!n308) & (!n376)) + ((!n121) & (n241) & (!n308) & (n376)) + ((!n121) & (n241) & (n308) & (n376)) + ((n121) & (n241) & (!n308) & (!n376)) + ((n121) & (n241) & (!n308) & (n376)) + ((n121) & (n241) & (n308) & (n376)));
	assign n201 = (((n203) & (n204) & (!n324) & (!n367)) + ((n203) & (n204) & (!n324) & (n367)) + ((n203) & (n204) & (n324) & (!n367)));
	assign n206 = (((!i_32_) & (!i_28_) & (n134)) + ((!i_32_) & (i_28_) & (!n134)) + ((!i_32_) & (i_28_) & (n134)) + ((i_32_) & (!i_28_) & (!n134)) + ((i_32_) & (!i_28_) & (n134)) + ((i_32_) & (i_28_) & (!n134)) + ((i_32_) & (i_28_) & (n134)));
	assign n205 = (((!n201) & (n206) & (!n394)) + ((n201) & (n206) & (!n394)) + ((n201) & (n206) & (n394)));
	assign n211 = (((!i_31_) & (!n253)) + ((!i_31_) & (n253)) + ((i_31_) & (!n253)));
	assign n207 = (((!i_30_) & (!i_32_) & (n211) & (!n253)) + ((!i_30_) & (!i_32_) & (n211) & (n253)) + ((!i_30_) & (i_32_) & (n211) & (!n253)) + ((i_30_) & (!i_32_) & (n211) & (!n253)) + ((i_30_) & (i_32_) & (n211) & (!n253)));
	assign n213 = (((!i_23_) & (!n957)) + ((i_23_) & (!n957)) + ((i_23_) & (n957)));
	assign n215 = (((!i_27_) & (n960)) + ((i_27_) & (!n960)) + ((i_27_) & (n960)));
	assign n216 = (((!i_14_) & (!n734)) + ((!i_14_) & (n734)) + ((i_14_) & (n734)));
	assign n212 = (((!n213) & (!n215) & (n216) & (!n363)) + ((!n213) & (n215) & (!n216) & (!n363)) + ((!n213) & (n215) & (n216) & (!n363)) + ((n213) & (!n215) & (n216) & (!n363)) + ((n213) & (!n215) & (n216) & (n363)) + ((n213) & (n215) & (!n216) & (!n363)) + ((n213) & (n215) & (!n216) & (n363)) + ((n213) & (n215) & (n216) & (!n363)) + ((n213) & (n215) & (n216) & (n363)));
	assign n219 = (((!i_20_) & (!n681) & (!n874) & (!n954)) + ((!i_20_) & (!n681) & (!n874) & (n954)) + ((!i_20_) & (!n681) & (n874) & (!n954)) + ((!i_20_) & (!n681) & (n874) & (n954)) + ((!i_20_) & (n681) & (!n874) & (!n954)) + ((!i_20_) & (n681) & (!n874) & (n954)) + ((!i_20_) & (n681) & (n874) & (!n954)) + ((!i_20_) & (n681) & (n874) & (n954)) + ((i_20_) & (!n681) & (!n874) & (!n954)) + ((i_20_) & (!n681) & (!n874) & (n954)) + ((i_20_) & (!n681) & (n874) & (!n954)) + ((i_20_) & (!n681) & (n874) & (n954)) + ((i_20_) & (n681) & (!n874) & (n954)) + ((i_20_) & (n681) & (n874) & (!n954)) + ((i_20_) & (n681) & (n874) & (n954)));
	assign n217 = (((!n212) & (n219) & (!n253) & (!n673)) + ((!n212) & (n219) & (!n253) & (n673)) + ((!n212) & (n219) & (n253) & (!n673)) + ((n212) & (n219) & (!n253) & (!n673)) + ((n212) & (n219) & (!n253) & (n673)) + ((n212) & (n219) & (n253) & (!n673)) + ((n212) & (n219) & (n253) & (n673)));
	assign n222 = (((!i_22_) & (!n256)) + ((i_22_) & (!n256)) + ((i_22_) & (n256)));
	assign n221 = (((!i_3_) & (!n22) & (n222)) + ((i_3_) & (!n22) & (!n222)) + ((i_3_) & (!n22) & (n222)));
	assign n224 = (((!i_7_) & (n177) & (!i_8_) & (n132)) + ((!i_7_) & (n177) & (i_8_) & (!n132)) + ((!i_7_) & (n177) & (i_8_) & (n132)) + ((i_7_) & (!n177) & (!i_8_) & (n132)) + ((i_7_) & (!n177) & (i_8_) & (!n132)) + ((i_7_) & (!n177) & (i_8_) & (n132)) + ((i_7_) & (n177) & (!i_8_) & (n132)) + ((i_7_) & (n177) & (i_8_) & (!n132)) + ((i_7_) & (n177) & (i_8_) & (n132)));
	assign n225 = (((!n224) & (n39) & (!n53) & (n221)) + ((!n224) & (n39) & (n53) & (!n221)) + ((!n224) & (n39) & (n53) & (n221)) + ((n224) & (!n39) & (!n53) & (n221)) + ((n224) & (!n39) & (n53) & (!n221)) + ((n224) & (!n39) & (n53) & (n221)) + ((n224) & (n39) & (!n53) & (n221)) + ((n224) & (n39) & (n53) & (!n221)) + ((n224) & (n39) & (n53) & (n221)));
	assign n227 = (((!i_22_) & (!n199)));
	assign n229 = (((!i_7_) & (!i_8_)));
	assign n226 = (((!n136) & (n227) & (n229)));
	assign n232 = (((i_12_) & (n23)));
	assign n230 = (((!i_11_) & (!n224) & (n226) & (n232)) + ((!i_11_) & (n224) & (n226) & (n232)) + ((i_11_) & (!n224) & (!n226) & (n232)) + ((i_11_) & (!n224) & (n226) & (n232)) + ((i_11_) & (n224) & (n226) & (n232)));
	assign n236 = (((!i_34_) & (!n995)) + ((!i_34_) & (n995)) + ((i_34_) & (n995)));
	assign n234 = (((!i_30_) & (!i_32_)));
	assign n233 = (((!i_28_) & (!i_34_) & (n236) & (!n234)) + ((!i_28_) & (!i_34_) & (n236) & (n234)) + ((!i_28_) & (i_34_) & (n236) & (n234)) + ((i_28_) & (!i_34_) & (n236) & (!n234)) + ((i_28_) & (!i_34_) & (n236) & (n234)) + ((i_28_) & (i_34_) & (n236) & (!n234)) + ((i_28_) & (i_34_) & (n236) & (n234)));
	assign n239 = (((!i_22_) & (!n234) & (!n233) & (!n356)) + ((!i_22_) & (!n234) & (n233) & (!n356)) + ((!i_22_) & (n234) & (!n233) & (!n356)) + ((!i_22_) & (n234) & (!n233) & (n356)) + ((!i_22_) & (n234) & (n233) & (!n356)) + ((!i_22_) & (n234) & (n233) & (n356)) + ((i_22_) & (!n234) & (n233) & (!n356)) + ((i_22_) & (n234) & (n233) & (!n356)) + ((i_22_) & (n234) & (n233) & (n356)));
	assign n238 = (((!i_29_) & (n724)) + ((i_29_) & (!n724)) + ((i_29_) & (n724)));
	assign n237 = (((n239) & (!i_28_) & (n238)) + ((n239) & (i_28_) & (!n238)) + ((n239) & (i_28_) & (n238)));
	assign n241 = (((!i_29_) & (n970)) + ((i_29_) & (!n970)) + ((i_29_) & (n970)));
	assign n240 = (((!i_25_) & (!i_28_) & (n241) & (!n367)) + ((!i_25_) & (i_28_) & (!n241) & (!n367)) + ((!i_25_) & (i_28_) & (n241) & (!n367)) + ((i_25_) & (!i_28_) & (n241) & (!n367)) + ((i_25_) & (!i_28_) & (n241) & (n367)) + ((i_25_) & (i_28_) & (!n241) & (!n367)) + ((i_25_) & (i_28_) & (!n241) & (n367)) + ((i_25_) & (i_28_) & (n241) & (!n367)) + ((i_25_) & (i_28_) & (n241) & (n367)));
	assign n243 = (((!i_31_) & (n974)) + ((i_31_) & (!n974)) + ((i_31_) & (n974)));
	assign n242 = (((!n92) & (n174) & (!i_8_) & (n243)) + ((!n92) & (n174) & (i_8_) & (!n243)) + ((!n92) & (n174) & (i_8_) & (n243)) + ((n92) & (!n174) & (!i_8_) & (n243)) + ((n92) & (!n174) & (i_8_) & (!n243)) + ((n92) & (!n174) & (i_8_) & (n243)) + ((n92) & (n174) & (!i_8_) & (n243)) + ((n92) & (n174) & (i_8_) & (!n243)) + ((n92) & (n174) & (i_8_) & (n243)));
	assign n246 = (((i_33_) & (n253)));
	assign n245 = (((i_33_) & (i_34_)));
	assign n244 = (((i_14_) & (!i_24_) & (!n246) & (n245)) + ((i_14_) & (!i_24_) & (n246) & (!n245)) + ((i_14_) & (!i_24_) & (n246) & (n245)) + ((i_14_) & (i_24_) & (n246) & (!n245)) + ((i_14_) & (i_24_) & (n246) & (n245)));
	assign n248 = (((n1012) & (n96)));
	assign n249 = (((!i_2_) & (!n229)) + ((i_2_) & (!n229)) + ((i_2_) & (n229)));
	assign n247 = (((!i_32_) & (n248) & (!i_30_) & (n249)) + ((!i_32_) & (n248) & (i_30_) & (!n249)) + ((!i_32_) & (n248) & (i_30_) & (n249)) + ((i_32_) & (!n248) & (!i_30_) & (n249)) + ((i_32_) & (!n248) & (i_30_) & (!n249)) + ((i_32_) & (!n248) & (i_30_) & (n249)) + ((i_32_) & (n248) & (!i_30_) & (n249)) + ((i_32_) & (n248) & (i_30_) & (!n249)) + ((i_32_) & (n248) & (i_30_) & (n249)));
	assign n250 = (((i_22_) & (!n207) & (!n213) & (n244)) + ((i_22_) & (!n207) & (n213) & (!n244)) + ((i_22_) & (!n207) & (n213) & (n244)) + ((i_22_) & (n207) & (!n213) & (n244)) + ((i_22_) & (n207) & (n213) & (n244)));
	assign n253 = (((!i_34_) & (i_35_)));
	assign n252 = (((!n29) & (!n253) & (!n290) & (!n1097)) + ((!n29) & (n253) & (!n290) & (!n1097)) + ((n29) & (!n253) & (!n290) & (!n1097)) + ((n29) & (n253) & (!n290) & (!n1097)) + ((n29) & (n253) & (!n290) & (n1097)));
	assign n256 = (((!i_13_) & (i_19_)));
	assign n255 = (((!n44) & (!n182) & (n256)) + ((n44) & (!n182) & (!n256)) + ((n44) & (!n182) & (n256)));
	assign n258 = (((!i_24_) & (!n23) & (!n74) & (n255)) + ((!i_24_) & (!n23) & (n74) & (n255)) + ((!i_24_) & (n23) & (!n74) & (!n255)) + ((!i_24_) & (n23) & (!n74) & (n255)) + ((!i_24_) & (n23) & (n74) & (n255)));
	assign n261 = (((!i_13_) & (n964)) + ((i_13_) & (!n964)) + ((i_13_) & (n964)));
	assign n260 = (((!i_18_) & (!n199) & (!n258) & (!n261)) + ((!i_18_) & (!n199) & (!n258) & (n261)) + ((!i_18_) & (n199) & (!n258) & (!n261)) + ((!i_18_) & (n199) & (!n258) & (n261)) + ((i_18_) & (!n199) & (!n258) & (n261)) + ((i_18_) & (n199) & (!n258) & (!n261)) + ((i_18_) & (n199) & (!n258) & (n261)));
	assign n263 = (((!i_18_) & (n39) & (!n44)) + ((!i_18_) & (n39) & (n44)) + ((i_18_) & (n39) & (!n44)));
	assign n266 = (((!n74) & (!n188) & (!n232) & (n263)) + ((!n74) & (n188) & (!n232) & (!n263)) + ((!n74) & (n188) & (!n232) & (n263)) + ((n74) & (!n188) & (!n232) & (n263)) + ((n74) & (!n188) & (n232) & (n263)) + ((n74) & (n188) & (!n232) & (!n263)) + ((n74) & (n188) & (!n232) & (n263)) + ((n74) & (n188) & (n232) & (!n263)) + ((n74) & (n188) & (n232) & (n263)));
	assign n265 = (((!i_12_) & (!n964)) + ((!i_12_) & (n964)) + ((i_12_) & (n964)));
	assign n264 = (((n266) & (!n39) & (n265)) + ((n266) & (n39) & (!n265)) + ((n266) & (n39) & (n265)));
	assign n268 = (((i_12_) & (n44)));
	assign n267 = (((i_18_) & (!i_22_) & (n268)));
	assign n269 = (((!i_8_) & (i_12_) & (!i_13_) & (n227) & (!n987)));
	assign n272 = (((!n90) & (n133) & (!n134) & (!n800)) + ((!n90) & (n133) & (n134) & (!n800)) + ((!n90) & (n133) & (n134) & (n800)) + ((n90) & (!n133) & (!n134) & (!n800)) + ((n90) & (!n133) & (n134) & (!n800)) + ((n90) & (!n133) & (n134) & (n800)) + ((n90) & (n133) & (!n134) & (!n800)) + ((n90) & (n133) & (n134) & (!n800)) + ((n90) & (n133) & (n134) & (n800)));
	assign n273 = (((!i_7_) & (n177) & (!n49) & (n221)) + ((!i_7_) & (n177) & (n49) & (!n221)) + ((!i_7_) & (n177) & (n49) & (n221)) + ((i_7_) & (!n177) & (!n49) & (n221)) + ((i_7_) & (!n177) & (n49) & (!n221)) + ((i_7_) & (!n177) & (n49) & (n221)) + ((i_7_) & (n177) & (!n49) & (n221)) + ((i_7_) & (n177) & (n49) & (!n221)) + ((i_7_) & (n177) & (n49) & (n221)));
	assign n274 = (((!i_2_) & (!i_10_) & (!i_12_) & (!n272)) + ((!i_2_) & (!i_10_) & (i_12_) & (!n272)) + ((i_2_) & (!i_10_) & (i_12_) & (!n272)));
	assign n282 = (((!i_3_) & (i_11_)));
	assign n279 = (((i_12_) & (!i_13_) & (!i_22_)));
	assign n278 = (((!n49) & (n282) & (!n279) & (!n1088)) + ((!n49) & (n282) & (n279) & (!n1088)) + ((!n49) & (n282) & (n279) & (n1088)) + ((n49) & (n282) & (!n279) & (!n1088)) + ((n49) & (n282) & (n279) & (!n1088)));
	assign n283 = (((!i_8_) & (!n19) & (n67) & (!n70)) + ((!i_8_) & (!n19) & (n67) & (n70)) + ((!i_8_) & (n19) & (n67) & (n70)) + ((i_8_) & (!n19) & (!n67) & (!n70)) + ((i_8_) & (!n19) & (!n67) & (n70)) + ((i_8_) & (!n19) & (n67) & (!n70)) + ((i_8_) & (!n19) & (n67) & (n70)) + ((i_8_) & (n19) & (!n67) & (n70)) + ((i_8_) & (n19) & (n67) & (n70)));
	assign n284 = (((!i_24_) & (!n66) & (!n69) & (!n240)));
	assign n288 = (((!i_24_) & (!i_25_)));
	assign n287 = (((!i_7_) & (!i_32_) & (n11) & (n288)));
	assign n290 = (((!i_31_) & (n234)));
	assign n289 = (((!i_22_) & (!i_23_) & (!n29) & (!n290)) + ((!i_22_) & (!i_23_) & (!n29) & (n290)) + ((!i_22_) & (!i_23_) & (n29) & (n290)) + ((!i_22_) & (i_23_) & (!n29) & (!n290)) + ((!i_22_) & (i_23_) & (!n29) & (n290)) + ((!i_22_) & (i_23_) & (n29) & (n290)) + ((i_22_) & (!i_23_) & (!n29) & (!n290)) + ((i_22_) & (!i_23_) & (!n29) & (n290)) + ((i_22_) & (!i_23_) & (n29) & (n290)));
	assign n293 = (((!i_38_) & (!n17) & (!n152) & (!n299)) + ((!i_38_) & (!n17) & (!n152) & (n299)) + ((!i_38_) & (!n17) & (n152) & (!n299)) + ((!i_38_) & (!n17) & (n152) & (n299)) + ((!i_38_) & (n17) & (!n152) & (!n299)) + ((!i_38_) & (n17) & (n152) & (!n299)) + ((i_38_) & (!n17) & (n152) & (!n299)) + ((i_38_) & (!n17) & (n152) & (n299)) + ((i_38_) & (n17) & (n152) & (!n299)));
	assign n299 = (((!i_31_) & (n394)));
	assign n296 = (((!i_29_) & (n299) & (!n1057)));
	assign n300 = (((!i_8_) & (!n11) & (!n288) & (!n299)) + ((!i_8_) & (!n11) & (!n288) & (n299)) + ((!i_8_) & (!n11) & (n288) & (!n299)) + ((!i_8_) & (!n11) & (n288) & (n299)) + ((!i_8_) & (n11) & (!n288) & (!n299)) + ((!i_8_) & (n11) & (!n288) & (n299)) + ((!i_8_) & (n11) & (n288) & (!n299)) + ((i_8_) & (!n11) & (!n288) & (!n299)) + ((i_8_) & (!n11) & (!n288) & (n299)) + ((i_8_) & (!n11) & (n288) & (!n299)) + ((i_8_) & (!n11) & (n288) & (n299)) + ((i_8_) & (n11) & (!n288) & (!n299)) + ((i_8_) & (n11) & (!n288) & (n299)) + ((i_8_) & (n11) & (n288) & (!n299)) + ((i_8_) & (n11) & (n288) & (n299)));
	assign n304 = (((!i_28_) & (n288)));
	assign n301 = (((!n190) & (!n296) & (n304) & (!n994)) + ((!n190) & (n296) & (n304) & (!n994)) + ((!n190) & (n296) & (n304) & (n994)) + ((n190) & (n296) & (n304) & (!n994)) + ((n190) & (n296) & (n304) & (n994)));
	assign n308 = (((!i_24_) & (n350)));
	assign n307 = (((!i_31_) & (n402) & (!n1057)));
	assign n306 = (((!i_30_) & (n402)));
	assign n305 = (((!n190) & (n308) & (!n307) & (n306)) + ((!n190) & (n308) & (n307) & (!n306)) + ((!n190) & (n308) & (n307) & (n306)) + ((n190) & (n308) & (n307) & (!n306)) + ((n190) & (n308) & (n307) & (n306)));
	assign n313 = (((!i_25_) & (n350)));
	assign n311 = (((n33) & (i_9_)));
	assign n309 = (((!n196) & (!n293) & (n313) & (!n311)) + ((!n196) & (!n293) & (n313) & (n311)) + ((!n196) & (n293) & (n313) & (n311)) + ((n196) & (!n293) & (n313) & (!n311)) + ((n196) & (!n293) & (n313) & (n311)));
	assign n315 = (((!i_29_) & (n995)) + ((i_29_) & (!n995)) + ((i_29_) & (n995)));
	assign n314 = (((!n35) & (!n315)) + ((!n35) & (n315)) + ((n35) & (n315)));
	assign n317 = (((i_38_) & (!n284) & (!n287) & (!n1081)) + ((i_38_) & (!n284) & (n287) & (!n1081)) + ((i_38_) & (!n284) & (n287) & (n1081)) + ((i_38_) & (n284) & (!n287) & (!n1081)) + ((i_38_) & (n284) & (!n287) & (n1081)) + ((i_38_) & (n284) & (n287) & (!n1081)) + ((i_38_) & (n284) & (n287) & (n1081)));
	assign n319 = (((!n86) & (!n139) & (n293) & (!n414)) + ((!n86) & (n139) & (n293) & (!n414)) + ((!n86) & (n139) & (n293) & (n414)) + ((n86) & (!n139) & (!n293) & (!n414)) + ((n86) & (!n139) & (n293) & (!n414)) + ((n86) & (n139) & (!n293) & (!n414)) + ((n86) & (n139) & (!n293) & (n414)) + ((n86) & (n139) & (n293) & (!n414)) + ((n86) & (n139) & (n293) & (n414)));
	assign n322 = (((!i_33_) & (i_38_)));
	assign n320 = (((!i_7_) & (!n163) & (n322)));
	assign n324 = (((!i_25_) & (!n163)));
	assign n323 = (((!i_32_) & (!n299) & (n320) & (!n324)) + ((!i_32_) & (!n299) & (n320) & (n324)) + ((!i_32_) & (n299) & (!n320) & (n324)) + ((!i_32_) & (n299) & (n320) & (!n324)) + ((!i_32_) & (n299) & (n320) & (n324)));
	assign n326 = (((!i_33_) & (!n299)) + ((i_33_) & (!n299)) + ((i_33_) & (n299)));
	assign n325 = (((!i_8_) & (!n163) & (!n323) & (n326)) + ((!i_8_) & (n163) & (!n323) & (!n326)) + ((!i_8_) & (n163) & (!n323) & (n326)) + ((i_8_) & (!n163) & (!n323) & (!n326)) + ((i_8_) & (!n163) & (!n323) & (n326)) + ((i_8_) & (n163) & (!n323) & (!n326)) + ((i_8_) & (n163) & (!n323) & (n326)));
	assign n328 = (((!i_25_) & (!n11) & (!n229) & (!n996)) + ((!i_25_) & (!n11) & (n229) & (!n996)) + ((!i_25_) & (n11) & (!n229) & (!n996)) + ((!i_25_) & (n11) & (n229) & (!n996)) + ((!i_25_) & (n11) & (n229) & (n996)));
	assign n331 = (((!i_32_) & (!n66) & (!n69) & (!n70)) + ((!i_32_) & (!n66) & (!n69) & (n70)) + ((!i_32_) & (n66) & (!n69) & (!n70)) + ((i_32_) & (!n66) & (!n69) & (!n70)) + ((i_32_) & (n66) & (!n69) & (!n70)));
	assign n335 = (((!n324) & (!n349) & (!n367) & (n1065)) + ((!n324) & (!n349) & (n367) & (n1065)) + ((!n324) & (n349) & (!n367) & (n1065)) + ((n324) & (!n349) & (!n367) & (n1065)) + ((n324) & (n349) & (!n367) & (n1065)));
	assign n336 = (((!n308) & (!n376) & (n1066)) + ((!n308) & (n376) & (n1066)) + ((n308) & (n376) & (n1066)));
	assign n334 = (((!i_32_) & (!n253)) + ((i_32_) & (!n253)) + ((i_32_) & (n253)));
	assign n332 = (((!n313) & (n335) & (n336) & (!n334)) + ((!n313) & (n335) & (n336) & (n334)) + ((n313) & (n335) & (n336) & (n334)));
	assign n337 = (((!i_7_) & (!n95) & (!n195) & (!n234)) + ((!i_7_) & (!n95) & (!n195) & (n234)) + ((!i_7_) & (n95) & (!n195) & (n234)) + ((i_7_) & (!n95) & (!n195) & (!n234)) + ((i_7_) & (!n95) & (!n195) & (n234)));
	assign n341 = (((!n66) & (!n350) & (!n716)) + ((!n66) & (!n350) & (n716)) + ((!n66) & (n350) & (n716)) + ((n66) & (!n350) & (!n716)) + ((n66) & (!n350) & (n716)) + ((n66) & (n350) & (!n716)) + ((n66) & (n350) & (n716)));
	assign n340 = (((!i_34_) & (!i_33_) & (i_29_)) + ((!i_34_) & (i_33_) & (!i_29_)) + ((!i_34_) & (i_33_) & (i_29_)) + ((i_34_) & (!i_33_) & (!i_29_)) + ((i_34_) & (!i_33_) & (i_29_)) + ((i_34_) & (i_33_) & (!i_29_)) + ((i_34_) & (i_33_) & (i_29_)));
	assign n339 = (((n341) & (!i_28_) & (!n70) & (n340)) + ((n341) & (!i_28_) & (n70) & (!n340)) + ((n341) & (!i_28_) & (n70) & (n340)) + ((n341) & (i_28_) & (!n70) & (!n340)) + ((n341) & (i_28_) & (!n70) & (n340)) + ((n341) & (i_28_) & (n70) & (!n340)) + ((n341) & (i_28_) & (n70) & (n340)));
	assign n342 = (((!n101) & (!n121) & (!n304) & (!n832)) + ((!n101) & (!n121) & (!n304) & (n832)) + ((!n101) & (!n121) & (n304) & (!n832)) + ((n101) & (!n121) & (!n304) & (!n832)) + ((n101) & (!n121) & (!n304) & (n832)) + ((n101) & (!n121) & (n304) & (!n832)) + ((n101) & (n121) & (!n304) & (!n832)) + ((n101) & (n121) & (!n304) & (n832)) + ((n101) & (n121) & (n304) & (!n832)));
	assign n345 = (((!i_33_) & (n978)) + ((i_33_) & (!n978)) + ((i_33_) & (n978)));
	assign n346 = (((!i_24_) & (i_28_)) + ((i_24_) & (!i_28_)) + ((i_24_) & (i_28_)));
	assign n347 = (((!i_33_) & (!n350)) + ((i_33_) & (!n350)) + ((i_33_) & (n350)));
	assign n344 = (((!n345) & (n346) & (!n163) & (n347)) + ((!n345) & (n346) & (n163) & (!n347)) + ((!n345) & (n346) & (n163) & (n347)) + ((n345) & (!n346) & (!n163) & (n347)) + ((n345) & (!n346) & (n163) & (!n347)) + ((n345) & (!n346) & (n163) & (n347)) + ((n345) & (n346) & (!n163) & (n347)) + ((n345) & (n346) & (n163) & (!n347)) + ((n345) & (n346) & (n163) & (n347)));
	assign n349 = (((!i_33_) & (n253)));
	assign n350 = (((!i_28_) & (!i_29_)));
	assign n348 = (((!n95) & (!n344) & (!n349) & (!n350)) + ((!n95) & (!n344) & (!n349) & (n350)) + ((!n95) & (!n344) & (n349) & (!n350)) + ((!n95) & (!n344) & (n349) & (n350)) + ((!n95) & (n344) & (n349) & (n350)));
	assign n352 = (((!n283) & (!n324) & (!n350) & (!n1062)) + ((!n283) & (!n324) & (n350) & (!n1062)) + ((!n283) & (n324) & (!n350) & (!n1062)) + ((!n283) & (n324) & (n350) & (!n1062)) + ((!n283) & (n324) & (n350) & (n1062)));
	assign n356 = (((n350) & (i_34_)));
	assign n355 = (((!n95) & (n288) & (!n356) & (!n1063)) + ((!n95) & (n288) & (n356) & (!n1063)) + ((!n95) & (n288) & (n356) & (n1063)) + ((n95) & (n288) & (!n356) & (!n1063)) + ((n95) & (n288) & (n356) & (!n1063)));
	assign n358 = (((n253) & (!n328) & (!n1067) & (!n1069)) + ((n253) & (!n328) & (!n1067) & (n1069)) + ((n253) & (!n328) & (n1067) & (!n1069)) + ((n253) & (n328) & (!n1067) & (!n1069)) + ((n253) & (n328) & (!n1067) & (n1069)) + ((n253) & (n328) & (n1067) & (!n1069)) + ((n253) & (n328) & (n1067) & (n1069)));
	assign n362 = (((!i_27_) & (n350)));
	assign n363 = (((n15) & (i_14_)));
	assign n364 = (((!i_16_) & (n833)));
	assign n361 = (((n362) & (n363) & (n364)));
	assign n367 = (((!i_32_) & (n350)));
	assign n365 = (((!n146) & (!n163) & (n367)));
	assign n368 = (((!n17) & (!n170) & (!n290) & (!n308)) + ((!n17) & (!n170) & (!n290) & (n308)) + ((!n17) & (!n170) & (n290) & (!n308)) + ((!n17) & (n170) & (!n290) & (!n308)) + ((!n17) & (n170) & (!n290) & (n308)) + ((!n17) & (n170) & (n290) & (!n308)) + ((n17) & (n170) & (!n290) & (!n308)) + ((n17) & (n170) & (!n290) & (n308)) + ((n17) & (n170) & (n290) & (!n308)));
	assign n371 = (((!i_5_) & (n961)) + ((i_5_) & (!n961)) + ((i_5_) & (n961)));
	assign n372 = (((!i_12_) & (i_6_)) + ((i_12_) & (!i_6_)) + ((i_12_) & (i_6_)));
	assign n373 = (((!i_5_) & (i_6_)) + ((i_5_) & (!i_6_)) + ((i_5_) & (i_6_)));
	assign n374 = (((!i_1_) & (n961)) + ((i_1_) & (!n961)) + ((i_1_) & (n961)));
	assign n370 = (((!n371) & (n372) & (!n373) & (n374)) + ((!n371) & (n372) & (n373) & (!n374)) + ((!n371) & (n372) & (n373) & (n374)) + ((n371) & (!n372) & (!n373) & (n374)) + ((n371) & (!n372) & (n373) & (!n374)) + ((n371) & (!n372) & (n373) & (n374)) + ((n371) & (n372) & (!n373) & (n374)) + ((n371) & (n372) & (n373) & (!n374)) + ((n371) & (n372) & (n373) & (n374)));
	assign n376 = (((!i_34_) & (!n970)) + ((!i_34_) & (n970)) + ((i_34_) & (n970)));
	assign n375 = (((!n190) & (!n311) & (!n324) & (!n376)) + ((!n190) & (!n311) & (!n324) & (n376)) + ((!n190) & (n311) & (!n324) & (n376)) + ((n190) & (!n311) & (!n324) & (!n376)) + ((n190) & (!n311) & (!n324) & (n376)) + ((n190) & (!n311) & (n324) & (!n376)) + ((n190) & (!n311) & (n324) & (n376)) + ((n190) & (n311) & (!n324) & (n376)) + ((n190) & (n311) & (n324) & (n376)));
	assign n377 = (((!i_29_) & (n140) & (!n192) & (!n311)) + ((!i_29_) & (n140) & (n192) & (!n311)) + ((!i_29_) & (n140) & (n192) & (n311)) + ((i_29_) & (!n140) & (!n192) & (!n311)) + ((i_29_) & (!n140) & (n192) & (!n311)) + ((i_29_) & (!n140) & (n192) & (n311)) + ((i_29_) & (n140) & (!n192) & (!n311)) + ((i_29_) & (n140) & (n192) & (!n311)) + ((i_29_) & (n140) & (n192) & (n311)));
	assign n378 = (((!i_24_) & (!n370) & (!n1045) & (!n1046)) + ((!i_24_) & (!n370) & (!n1045) & (n1046)) + ((!i_24_) & (!n370) & (n1045) & (!n1046)));
	assign n382 = (((!n86) & (n227) & (!n1258)) + ((!n86) & (n227) & (n1258)) + ((n86) & (n227) & (!n1258)));
	assign n385 = (((!n1047) & (!n1048) & (!n1049) & (!n1051)) + ((!n1047) & (!n1048) & (!n1049) & (n1051)) + ((!n1047) & (!n1048) & (n1049) & (!n1051)) + ((!n1047) & (n1048) & (!n1049) & (!n1051)) + ((!n1047) & (n1048) & (!n1049) & (n1051)) + ((!n1047) & (n1048) & (n1049) & (!n1051)) + ((n1047) & (!n1048) & (!n1049) & (!n1051)) + ((n1047) & (!n1048) & (!n1049) & (n1051)) + ((n1047) & (!n1048) & (n1049) & (!n1051)));
	assign n394 = (((!i_35_) & (i_38_)));
	assign n390 = (((n394) & (!n1053) & (!n1055) & (!n1058)) + ((n394) & (!n1053) & (!n1055) & (n1058)) + ((n394) & (!n1053) & (n1055) & (!n1058)) + ((n394) & (!n1053) & (n1055) & (n1058)) + ((n394) & (n1053) & (!n1055) & (!n1058)) + ((n394) & (n1053) & (!n1055) & (n1058)) + ((n394) & (n1053) & (n1055) & (!n1058)));
	assign n395 = (((!n185) & (!n283) & (!n307) & (n322)) + ((!n185) & (!n283) & (n307) & (!n322)) + ((!n185) & (!n283) & (n307) & (n322)) + ((!n185) & (n283) & (n307) & (!n322)) + ((!n185) & (n283) & (n307) & (n322)));
	assign n397 = (((!i_12_) & (!n181) & (!n256) & (n268)) + ((!i_12_) & (!n181) & (n256) & (n268)) + ((i_12_) & (!n181) & (!n256) & (n268)) + ((i_12_) & (!n181) & (n256) & (!n268)) + ((i_12_) & (!n181) & (n256) & (n268)));
	assign n402 = (((!i_33_) & (n394)));
	assign n399 = (((!n138) & (!n186) & (!n365) & (n402)) + ((!n138) & (!n186) & (n365) & (n402)) + ((!n138) & (n186) & (n365) & (n402)) + ((n138) & (!n186) & (n365) & (n402)) + ((n138) & (n186) & (n365) & (n402)));
	assign n404 = (((n362) & (!n608)));
	assign n403 = (((!n216) & (n245) & (!n361) & (n404)) + ((!n216) & (n245) & (n361) & (!n404)) + ((!n216) & (n245) & (n361) & (n404)) + ((n216) & (n245) & (n361) & (!n404)) + ((n216) & (n245) & (n361) & (n404)));
	assign n407 = (((n350) & (n290) & (n246)));
	assign n406 = (((i_14_) & (!n407) & (n121) & (i_33_)) + ((i_14_) & (n407) & (!n121) & (!i_33_)) + ((i_14_) & (n407) & (!n121) & (i_33_)) + ((i_14_) & (n407) & (n121) & (!i_33_)) + ((i_14_) & (n407) & (n121) & (i_33_)));
	assign n408 = (((i_9_) & (!n1089) & (!n1091) & (!n1093)) + ((i_9_) & (!n1089) & (!n1091) & (n1093)) + ((i_9_) & (!n1089) & (n1091) & (!n1093)) + ((i_9_) & (!n1089) & (n1091) & (n1093)) + ((i_9_) & (n1089) & (!n1091) & (!n1093)) + ((i_9_) & (n1089) & (!n1091) & (n1093)) + ((i_9_) & (n1089) & (n1091) & (!n1093)));
	assign n413 = (((i_10_) & (!n267) & (n282) & (n279)) + ((i_10_) & (n267) & (!n282) & (!n279)) + ((i_10_) & (n267) & (!n282) & (n279)) + ((i_10_) & (n267) & (n282) & (!n279)) + ((i_10_) & (n267) & (n282) & (n279)));
	assign n414 = (((!i_24_) & (n229)));
	assign n412 = (((!n136) & (!n269) & (n413) & (n414)) + ((!n136) & (n269) & (!n413) & (!n414)) + ((!n136) & (n269) & (!n413) & (n414)) + ((!n136) & (n269) & (n413) & (!n414)) + ((!n136) & (n269) & (n413) & (n414)));
	assign n415 = (((!i_28_) & (!n250) & (!n252) & (!n1263)) + ((!i_28_) & (!n250) & (n252) & (!n1263)) + ((!i_28_) & (!n250) & (n252) & (n1263)) + ((!i_28_) & (n250) & (!n252) & (!n1263)) + ((!i_28_) & (n250) & (!n252) & (n1263)) + ((!i_28_) & (n250) & (n252) & (!n1263)) + ((!i_28_) & (n250) & (n252) & (n1263)));
	assign n418 = (((i_10_) & (!i_12_) & (!n225) & (!n1102)) + ((i_10_) & (!i_12_) & (n225) & (!n1102)) + ((i_10_) & (i_12_) & (!n225) & (!n1102)) + ((i_10_) & (i_12_) & (!n225) & (n1102)) + ((i_10_) & (i_12_) & (n225) & (!n1102)));
	assign n421 = (((n48) & (!n127) & (!n997) & (!n1106)) + ((n48) & (!n127) & (!n997) & (n1106)) + ((n48) & (!n127) & (n997) & (!n1106)) + ((n48) & (n127) & (!n997) & (!n1106)) + ((n48) & (n127) & (n997) & (!n1106)));
	assign n425 = (((!n121) & (n213) & (!n234) & (!n1108)) + ((!n121) & (n213) & (n234) & (!n1108)) + ((n121) & (n213) & (!n234) & (!n1108)) + ((n121) & (n213) & (!n234) & (n1108)) + ((n121) & (n213) & (n234) & (!n1108)));
	assign n429 = (((!i_22_) & (n33)));
	assign n428 = (((!n85) & (!n371) & (!n429) & (!n1113)) + ((!n85) & (!n371) & (n429) & (!n1113)) + ((!n85) & (!n371) & (n429) & (n1113)) + ((n85) & (!n371) & (!n429) & (!n1113)) + ((n85) & (!n371) & (n429) & (!n1113)));
	assign n436 = (((!i_27_) & (!n179) & (!n390) & (!n531)) + ((!i_27_) & (!n179) & (!n390) & (n531)) + ((!i_27_) & (n179) & (!n390) & (!n531)) + ((!i_27_) & (n179) & (!n390) & (n531)) + ((i_27_) & (!n179) & (!n390) & (!n531)) + ((i_27_) & (n179) & (!n390) & (!n531)) + ((i_27_) & (n179) & (!n390) & (n531)));
	assign n437 = (((n1141) & (!n49) & (!n222) & (n969)) + ((n1141) & (!n49) & (n222) & (!n969)) + ((n1141) & (!n49) & (n222) & (n969)) + ((n1141) & (n49) & (!n222) & (!n969)) + ((n1141) & (n49) & (!n222) & (n969)) + ((n1141) & (n49) & (n222) & (!n969)) + ((n1141) & (n49) & (n222) & (n969)));
	assign n438 = (((!n35) & (!n234) & (!n356) & (n1139)) + ((!n35) & (!n234) & (n356) & (n1139)) + ((!n35) & (n234) & (!n356) & (n1139)) + ((!n35) & (n234) & (n356) & (n1139)) + ((n35) & (!n234) & (!n356) & (n1139)) + ((n35) & (n234) & (!n356) & (n1139)) + ((n35) & (n234) & (n356) & (n1139)));
	assign n439 = (((!n11) & (!n325) & (!n406) & (n1146)) + ((!n11) & (n325) & (!n406) & (n1146)) + ((n11) & (n325) & (!n406) & (n1146)));
	assign n440 = (((!n124) & (n368) & (!n399) & (n1143)) + ((n124) & (!n368) & (!n399) & (n1143)) + ((n124) & (n368) & (!n399) & (n1143)));
	assign n441 = (((!n418) & (!n421) & (n1149) & (n1152) & (n1153) & (n1157) & (n1159) & (n1160)));
	assign n433 = (((!n395) & (!n397) & (n436) & (n437) & (n438) & (n439) & (n440) & (n441)));
	assign n443 = (((!i_34_) & (!i_37_)) + ((!i_34_) & (i_37_)) + ((i_34_) & (!i_37_)));
	assign n444 = (((!i_29_) & (n649)) + ((i_29_) & (!n649)) + ((i_29_) & (n649)));
	assign n446 = (((!i_37_) & (!n253)) + ((!i_37_) & (n253)) + ((i_37_) & (!n253)));
	assign n442 = (((!n362) & (!n443) & (n444) & (!n446)) + ((!n362) & (!n443) & (n444) & (n446)) + ((!n362) & (n443) & (!n444) & (!n446)) + ((!n362) & (n443) & (!n444) & (n446)) + ((!n362) & (n443) & (n444) & (!n446)) + ((!n362) & (n443) & (n444) & (n446)) + ((n362) & (!n443) & (n444) & (n446)) + ((n362) & (n443) & (!n444) & (n446)) + ((n362) & (n443) & (n444) & (n446)));
	assign n449 = (((!i_29_) & (!n543) & (!n664)) + ((!i_29_) & (!n543) & (n664)) + ((!i_29_) & (n543) & (n664)) + ((i_29_) & (!n543) & (!n664)) + ((i_29_) & (!n543) & (n664)) + ((i_29_) & (n543) & (!n664)) + ((i_29_) & (n543) & (n664)));
	assign n448 = (((!i_34_) & (!n543)) + ((!i_34_) & (n543)) + ((i_34_) & (!n543)));
	assign n447 = (((!n362) & (n449) & (!n448)) + ((!n362) & (n449) & (n448)) + ((n362) & (n449) & (n448)));
	assign n451 = (((!i_37_) & (!n362) & (!n832)) + ((!i_37_) & (!n362) & (n832)) + ((!i_37_) & (n362) & (!n832)) + ((!i_37_) & (n362) & (n832)) + ((i_37_) & (!n362) & (!n832)) + ((i_37_) & (!n362) & (n832)) + ((i_37_) & (n362) & (!n832)));
	assign n450 = (((n451) & (!i_32_) & (n449)) + ((n451) & (i_32_) & (!n449)) + ((n451) & (i_32_) & (n449)));
	assign n455 = (((!n371) & (!n453) & (n1020)) + ((!n371) & (n453) & (!n1020)) + ((!n371) & (n453) & (n1020)) + ((n371) & (!n453) & (!n1020)) + ((n371) & (!n453) & (n1020)) + ((n371) & (n453) & (!n1020)) + ((n371) & (n453) & (n1020)));
	assign n453 = (((!i_17_) & (n735)) + ((i_17_) & (!n735)) + ((i_17_) & (n735)));
	assign n454 = (((!i_10_) & (n989)) + ((i_10_) & (!n989)) + ((i_10_) & (n989)));
	assign n452 = (((n455) & (!n371) & (!n453) & (n454)) + ((n455) & (!n371) & (n453) & (!n454)) + ((n455) & (!n371) & (n453) & (n454)) + ((n455) & (n371) & (!n453) & (!n454)) + ((n455) & (n371) & (!n453) & (n454)) + ((n455) & (n371) & (n453) & (!n454)) + ((n455) & (n371) & (n453) & (n454)));
	assign n459 = (((!n1015) & (!n454) & (!n522) & (n501)) + ((!n1015) & (!n454) & (n522) & (!n501)) + ((!n1015) & (!n454) & (n522) & (n501)) + ((!n1015) & (n454) & (!n522) & (!n501)) + ((!n1015) & (n454) & (!n522) & (n501)) + ((!n1015) & (n454) & (n522) & (!n501)) + ((!n1015) & (n454) & (n522) & (n501)) + ((n1015) & (!n454) & (!n522) & (!n501)) + ((n1015) & (!n454) & (!n522) & (n501)) + ((n1015) & (!n454) & (n522) & (!n501)) + ((n1015) & (!n454) & (n522) & (n501)) + ((n1015) & (n454) & (!n522) & (!n501)) + ((n1015) & (n454) & (!n522) & (n501)) + ((n1015) & (n454) & (n522) & (!n501)) + ((n1015) & (n454) & (n522) & (n501)));
	assign n457 = (((!i_37_) & (!n595) & (!n622)) + ((!i_37_) & (!n595) & (n622)) + ((!i_37_) & (n595) & (!n622)) + ((!i_37_) & (n595) & (n622)) + ((i_37_) & (!n595) & (n622)) + ((i_37_) & (n595) & (!n622)) + ((i_37_) & (n595) & (n622)));
	assign n458 = (((!n543) & (!n1015) & (!n1114)) + ((!n543) & (!n1015) & (n1114)) + ((!n543) & (n1015) & (!n1114)) + ((!n543) & (n1015) & (n1114)) + ((n543) & (!n1015) & (n1114)) + ((n543) & (n1015) & (!n1114)) + ((n543) & (n1015) & (n1114)));
	assign n456 = (((n459) & (!n453) & (n457) & (n458)) + ((n459) & (n453) & (!n457) & (!n458)) + ((n459) & (n453) & (!n457) & (n458)) + ((n459) & (n453) & (n457) & (!n458)) + ((n459) & (n453) & (n457) & (n458)));
	assign n462 = (((!n494) & (!n992) & (!n1015)) + ((!n494) & (!n992) & (n1015)) + ((!n494) & (n992) & (!n1015)) + ((!n494) & (n992) & (n1015)) + ((n494) & (!n992) & (n1015)) + ((n494) & (n992) & (!n1015)) + ((n494) & (n992) & (n1015)));
	assign n461 = (((!i_7_) & (!i_0_) & (n1005)) + ((!i_7_) & (i_0_) & (!n1005)) + ((!i_7_) & (i_0_) & (n1005)) + ((i_7_) & (!i_0_) & (!n1005)) + ((i_7_) & (!i_0_) & (n1005)) + ((i_7_) & (i_0_) & (!n1005)) + ((i_7_) & (i_0_) & (n1005)));
	assign n460 = (((n462) & (!i_12_) & (n461)) + ((n462) & (i_12_) & (!n461)) + ((n462) & (i_12_) & (n461)));
	assign n467 = (((!i_23_) & (!n163)));
	assign n463 = (((!n460) & (n467) & (!n629) & (!n1194)) + ((!n460) & (n467) & (!n629) & (n1194)) + ((!n460) & (n467) & (n629) & (!n1194)) + ((n460) & (n467) & (!n629) & (!n1194)) + ((n460) & (n467) & (n629) & (!n1194)));
	assign n471 = (((!n639) & (!n1009) & (n587)) + ((!n639) & (n1009) & (!n587)) + ((!n639) & (n1009) & (n587)) + ((n639) & (!n1009) & (!n587)) + ((n639) & (!n1009) & (n587)) + ((n639) & (n1009) & (!n587)) + ((n639) & (n1009) & (n587)));
	assign n469 = (((!i_11_) & (n735)) + ((i_11_) & (!n735)) + ((i_11_) & (n735)));
	assign n470 = (((!n81) & (!n1015) & (n746)) + ((!n81) & (n1015) & (!n746)) + ((!n81) & (n1015) & (n746)) + ((n81) & (!n1015) & (!n746)) + ((n81) & (!n1015) & (n746)) + ((n81) & (n1015) & (!n746)) + ((n81) & (n1015) & (n746)));
	assign n468 = (((!n463) & (n471) & (!n469) & (n470)) + ((!n463) & (n471) & (n469) & (!n470)) + ((!n463) & (n471) & (n469) & (n470)));
	assign n474 = (((!i_14_) & (!n543)) + ((i_14_) & (!n543)) + ((i_14_) & (n543)));
	assign n473 = (((!i_21_) & (!n11) & (!n474) & (!n692)) + ((!i_21_) & (!n11) & (!n474) & (n692)) + ((!i_21_) & (!n11) & (n474) & (!n692)) + ((!i_21_) & (!n11) & (n474) & (n692)) + ((!i_21_) & (n11) & (n474) & (!n692)) + ((!i_21_) & (n11) & (n474) & (n692)) + ((i_21_) & (!n11) & (!n474) & (!n692)) + ((i_21_) & (!n11) & (n474) & (!n692)) + ((i_21_) & (n11) & (n474) & (!n692)));
	assign n479 = (((n953) & (n453)));
	assign n477 = (((!i_33_) & (n479) & (!n688)) + ((i_33_) & (n479) & (!n688)) + ((i_33_) & (n479) & (n688)));
	assign n482 = (((!n66) & (n763)) + ((n66) & (!n763)) + ((n66) & (n763)));
	assign n481 = (((!i_10_) & (n735)) + ((i_10_) & (!n735)) + ((i_10_) & (n735)));
	assign n480 = (((n482) & (!n66) & (n481)) + ((n482) & (n66) & (!n481)) + ((n482) & (n66) & (n481)));
	assign n485 = (((!i_31_) & (!n11) & (!n477) & (!n572)) + ((!i_31_) & (!n11) & (!n477) & (n572)) + ((!i_31_) & (!n11) & (n477) & (!n572)) + ((!i_31_) & (!n11) & (n477) & (n572)) + ((!i_31_) & (n11) & (!n477) & (!n572)) + ((!i_31_) & (n11) & (!n477) & (n572)) + ((!i_31_) & (n11) & (n477) & (!n572)) + ((!i_31_) & (n11) & (n477) & (n572)) + ((i_31_) & (!n11) & (!n477) & (!n572)) + ((i_31_) & (!n11) & (!n477) & (n572)) + ((i_31_) & (!n11) & (n477) & (!n572)) + ((i_31_) & (!n11) & (n477) & (n572)) + ((i_31_) & (n11) & (!n477) & (n572)) + ((i_31_) & (n11) & (n477) & (!n572)) + ((i_31_) & (n11) & (n477) & (n572)));
	assign n483 = (((!n404) & (!n480) & (n485)) + ((!n404) & (n480) & (n485)) + ((n404) & (n480) & (n485)));
	assign n487 = (((!i_29_) & (!n456) & (!n664) & (!n1027)) + ((!i_29_) & (!n456) & (!n664) & (n1027)) + ((!i_29_) & (!n456) & (n664) & (!n1027)) + ((!i_29_) & (!n456) & (n664) & (n1027)) + ((!i_29_) & (n456) & (!n664) & (!n1027)) + ((!i_29_) & (n456) & (!n664) & (n1027)) + ((!i_29_) & (n456) & (n664) & (!n1027)) + ((!i_29_) & (n456) & (n664) & (n1027)) + ((i_29_) & (!n456) & (!n664) & (n1027)) + ((i_29_) & (!n456) & (n664) & (!n1027)) + ((i_29_) & (!n456) & (n664) & (n1027)) + ((i_29_) & (n456) & (!n664) & (!n1027)) + ((i_29_) & (n456) & (!n664) & (n1027)) + ((i_29_) & (n456) & (n664) & (!n1027)) + ((i_29_) & (n456) & (n664) & (n1027)));
	assign n488 = (((!n884) & (!n561) & (!n1023) & (i_29_)) + ((!n884) & (!n561) & (n1023) & (!i_29_)) + ((!n884) & (!n561) & (n1023) & (i_29_)) + ((!n884) & (n561) & (!n1023) & (!i_29_)) + ((!n884) & (n561) & (!n1023) & (i_29_)) + ((!n884) & (n561) & (n1023) & (!i_29_)) + ((!n884) & (n561) & (n1023) & (i_29_)) + ((n884) & (!n561) & (!n1023) & (!i_29_)) + ((n884) & (!n561) & (!n1023) & (i_29_)) + ((n884) & (!n561) & (n1023) & (!i_29_)) + ((n884) & (!n561) & (n1023) & (i_29_)) + ((n884) & (n561) & (!n1023) & (!i_29_)) + ((n884) & (n561) & (!n1023) & (i_29_)) + ((n884) & (n561) & (n1023) & (!i_29_)) + ((n884) & (n561) & (n1023) & (i_29_)));
	assign n489 = (((!i_37_) & (!n443) & (!n468) & (n483)) + ((!i_37_) & (!n443) & (n468) & (n483)) + ((!i_37_) & (n443) & (!n468) & (!n483)) + ((!i_37_) & (n443) & (!n468) & (n483)) + ((!i_37_) & (n443) & (n468) & (!n483)) + ((!i_37_) & (n443) & (n468) & (n483)) + ((i_37_) & (!n443) & (n468) & (n483)) + ((i_37_) & (n443) & (n468) & (!n483)) + ((i_37_) & (n443) & (n468) & (n483)));
	assign n490 = (((n1196) & (!i_31_) & (!n473) & (n684)) + ((n1196) & (!i_31_) & (n473) & (!n684)) + ((n1196) & (!i_31_) & (n473) & (n684)) + ((n1196) & (i_31_) & (!n473) & (!n684)) + ((n1196) & (i_31_) & (!n473) & (n684)) + ((n1196) & (i_31_) & (n473) & (!n684)) + ((n1196) & (i_31_) & (n473) & (n684)));
	assign n486 = (((n487) & (n488) & (n489) & (n490)));
	assign n494 = (((!i_27_) & (n531)));
	assign n495 = (((n833) & (i_22_)));
	assign n491 = (((!n479) & (n494) & (n495) & (!n1011)) + ((!n479) & (n494) & (n495) & (n1011)) + ((n479) & (n494) & (n495) & (!n1011)));
	assign n497 = (((!i_33_) & (!n685)) + ((!i_33_) & (n685)) + ((i_33_) & (n685)));
	assign n498 = (((!i_25_) & (!n833)) + ((!i_25_) & (n833)) + ((i_25_) & (!n833)));
	assign n496 = (((!n11) & (!n491) & (!n497) & (!n498)) + ((!n11) & (!n491) & (!n497) & (n498)) + ((!n11) & (!n491) & (n497) & (!n498)) + ((!n11) & (!n491) & (n497) & (n498)) + ((n11) & (!n491) & (!n497) & (n498)) + ((n11) & (!n491) & (n497) & (!n498)) + ((n11) & (!n491) & (n497) & (n498)));
	assign n501 = (((!i_33_) & (!n543)) + ((i_33_) & (!n543)) + ((i_33_) & (n543)));
	assign n500 = (((n474) & (!i_13_) & (n501)) + ((n474) & (i_13_) & (!n501)) + ((n474) & (i_13_) & (n501)));
	assign n503 = (((n481) & (n763)));
	assign n505 = (((!i_10_) & (n734)) + ((i_10_) & (!n734)) + ((i_10_) & (n734)));
	assign n502 = (((!n501) & (!n503) & (n505) & (!n543)) + ((!n501) & (n503) & (n505) & (!n543)) + ((!n501) & (n503) & (n505) & (n543)) + ((n501) & (!n503) & (!n505) & (!n543)) + ((n501) & (!n503) & (n505) & (!n543)) + ((n501) & (n503) & (!n505) & (!n543)) + ((n501) & (n503) & (!n505) & (n543)) + ((n501) & (n503) & (n505) & (!n543)) + ((n501) & (n503) & (n505) & (n543)));
	assign n506 = (((!i_33_) & (!n457) & (!n609) & (!n620)) + ((!i_33_) & (!n457) & (!n609) & (n620)) + ((!i_33_) & (!n457) & (n609) & (!n620)) + ((i_33_) & (!n457) & (!n609) & (!n620)) + ((i_33_) & (!n457) & (n609) & (!n620)));
	assign n512 = (((!i_20_) & (!n1003)) + ((i_20_) & (!n1003)) + ((i_20_) & (n1003)));
	assign n513 = (((!i_20_) & (n960)) + ((i_20_) & (!n960)) + ((i_20_) & (n960)));
	assign n511 = (((!i_12_) & (n512) & (!i_16_) & (n513)) + ((!i_12_) & (n512) & (i_16_) & (!n513)) + ((!i_12_) & (n512) & (i_16_) & (n513)) + ((i_12_) & (!n512) & (!i_16_) & (n513)) + ((i_12_) & (!n512) & (i_16_) & (!n513)) + ((i_12_) & (!n512) & (i_16_) & (n513)) + ((i_12_) & (n512) & (!i_16_) & (n513)) + ((i_12_) & (n512) & (i_16_) & (!n513)) + ((i_12_) & (n512) & (i_16_) & (n513)));
	assign n516 = (((n1169) & (!n990) & (!n639) & (n1013)) + ((n1169) & (!n990) & (n639) & (!n1013)) + ((n1169) & (!n990) & (n639) & (n1013)) + ((n1169) & (n990) & (!n639) & (!n1013)) + ((n1169) & (n990) & (!n639) & (n1013)) + ((n1169) & (n990) & (n639) & (!n1013)) + ((n1169) & (n990) & (n639) & (n1013)));
	assign n515 = (((!i_19_) & (n960)) + ((i_19_) & (!n960)) + ((i_19_) & (n960)));
	assign n514 = (((n516) & (!n59) & (!n515) & (n469)) + ((n516) & (!n59) & (n515) & (!n469)) + ((n516) & (!n59) & (n515) & (n469)) + ((n516) & (n59) & (!n515) & (!n469)) + ((n516) & (n59) & (!n515) & (n469)) + ((n516) & (n59) & (n515) & (!n469)) + ((n516) & (n59) & (n515) & (n469)));
	assign n519 = (((!n990) & (!n640) & (n1013)) + ((!n990) & (n640) & (!n1013)) + ((!n990) & (n640) & (n1013)) + ((n990) & (!n640) & (!n1013)) + ((n990) & (!n640) & (n1013)) + ((n990) & (n640) & (!n1013)) + ((n990) & (n640) & (n1013)));
	assign n518 = (((!i_11_) & (n734)) + ((i_11_) & (!n734)) + ((i_11_) & (n734)));
	assign n517 = (((n519) & (!n59) & (!n515) & (n518)) + ((n519) & (!n59) & (n515) & (!n518)) + ((n519) & (!n59) & (n515) & (n518)) + ((n519) & (n59) & (!n515) & (!n518)) + ((n519) & (n59) & (!n515) & (n518)) + ((n519) & (n59) & (n515) & (!n518)) + ((n519) & (n59) & (n515) & (n518)));
	assign n520 = (((n503) & (!i_33_) & (n505)) + ((n503) & (i_33_) & (!n505)) + ((n503) & (i_33_) & (n505)));
	assign n522 = (((!i_17_) & (n734)) + ((i_17_) & (!n734)) + ((i_17_) & (n734)));
	assign n521 = (((!n453) & (!n501) & (n522) & (!n543)) + ((!n453) & (n501) & (!n522) & (!n543)) + ((!n453) & (n501) & (n522) & (!n543)) + ((n453) & (!n501) & (n522) & (!n543)) + ((n453) & (!n501) & (n522) & (n543)) + ((n453) & (n501) & (!n522) & (!n543)) + ((n453) & (n501) & (!n522) & (n543)) + ((n453) & (n501) & (n522) & (!n543)) + ((n453) & (n501) & (n522) & (n543)));
	assign n524 = (((n1192) & (!i_19_) & (!n991) & (n526)) + ((n1192) & (!i_19_) & (n991) & (!n526)) + ((n1192) & (!i_19_) & (n991) & (n526)) + ((n1192) & (i_19_) & (!n991) & (!n526)) + ((n1192) & (i_19_) & (!n991) & (n526)) + ((n1192) & (i_19_) & (n991) & (!n526)) + ((n1192) & (i_19_) & (n991) & (n526)));
	assign n523 = (((n524) & (!n500) & (!n372) & (n512)) + ((n524) & (!n500) & (n372) & (!n512)) + ((n524) & (!n500) & (n372) & (n512)) + ((n524) & (n500) & (!n372) & (!n512)) + ((n524) & (n500) & (!n372) & (n512)) + ((n524) & (n500) & (n372) & (!n512)) + ((n524) & (n500) & (n372) & (n512)));
	assign n526 = (((!i_23_) & (!i_20_) & (n521)) + ((!i_23_) & (i_20_) & (!n521)) + ((!i_23_) & (i_20_) & (n521)) + ((i_23_) & (!i_20_) & (!n521)) + ((i_23_) & (!i_20_) & (n521)) + ((i_23_) & (i_20_) & (!n521)) + ((i_23_) & (i_20_) & (n521)));
	assign n527 = (((!i_3_) & (!n1007)) + ((!i_3_) & (n1007)) + ((i_3_) & (n1007)));
	assign n528 = (((!i_9_) & (n373)) + ((i_9_) & (!n373)) + ((i_9_) & (n373)));
	assign n525 = (((!n526) & (!n527) & (!n528) & (i_18_)) + ((!n526) & (!n527) & (n528) & (!i_18_)) + ((!n526) & (!n527) & (n528) & (i_18_)) + ((!n526) & (n527) & (!n528) & (!i_18_)) + ((!n526) & (n527) & (!n528) & (i_18_)) + ((!n526) & (n527) & (n528) & (!i_18_)) + ((!n526) & (n527) & (n528) & (i_18_)) + ((n526) & (!n527) & (!n528) & (!i_18_)) + ((n526) & (!n527) & (!n528) & (i_18_)) + ((n526) & (!n527) & (n528) & (!i_18_)) + ((n526) & (!n527) & (n528) & (i_18_)) + ((n526) & (n527) & (!n528) & (!i_18_)) + ((n526) & (n527) & (!n528) & (i_18_)) + ((n526) & (n527) & (n528) & (!i_18_)) + ((n526) & (n527) & (n528) & (i_18_)));
	assign n531 = (((!i_28_) & (i_29_)));
	assign n529 = (((!n506) & (!n513) & (n531) & (!n1190)) + ((n506) & (!n513) & (n531) & (!n1190)) + ((n506) & (!n513) & (n531) & (n1190)));
	assign n534 = (((!i_13_) & (!n1014) & (n556)) + ((!i_13_) & (n1014) & (!n556)) + ((!i_13_) & (n1014) & (n556)) + ((i_13_) & (!n1014) & (!n556)) + ((i_13_) & (!n1014) & (n556)) + ((i_13_) & (n1014) & (!n556)) + ((i_13_) & (n1014) & (n556)));
	assign n533 = (((!n367) & (!n501) & (!n534)) + ((!n367) & (!n501) & (n534)) + ((!n367) & (n501) & (!n534)) + ((!n367) & (n501) & (n534)) + ((n367) & (!n501) & (n534)) + ((n367) & (n501) & (!n534)) + ((n367) & (n501) & (n534)));
	assign n539 = (((!i_32_) & (n531)));
	assign n535 = (((!n523) & (!n525) & (n539) & (!n1015)) + ((!n523) & (!n525) & (n539) & (n1015)) + ((!n523) & (n525) & (n539) & (!n1015)) + ((n523) & (!n525) & (n539) & (!n1015)) + ((n523) & (!n525) & (n539) & (n1015)));
	assign n543 = (((!i_35_) & (i_37_)));
	assign n540 = (((!n367) & (n543) & (!n704) & (!n1193)) + ((!n367) & (n543) & (n704) & (!n1193)) + ((n367) & (n543) & (!n704) & (!n1193)) + ((n367) & (n543) & (!n704) & (n1193)) + ((n367) & (n543) & (n704) & (!n1193)));
	assign n545 = (((n1163) & (!n984) & (!n640) & (n1013)) + ((n1163) & (!n984) & (n640) & (!n1013)) + ((n1163) & (!n984) & (n640) & (n1013)) + ((n1163) & (n984) & (!n640) & (!n1013)) + ((n1163) & (n984) & (!n640) & (n1013)) + ((n1163) & (n984) & (n640) & (!n1013)) + ((n1163) & (n984) & (n640) & (n1013)));
	assign n544 = (((n545) & (!n66) & (!n515) & (n518)) + ((n545) & (!n66) & (n515) & (!n518)) + ((n545) & (!n66) & (n515) & (n518)) + ((n545) & (n66) & (!n515) & (!n518)) + ((n545) & (n66) & (!n515) & (n518)) + ((n545) & (n66) & (n515) & (!n518)) + ((n545) & (n66) & (n515) & (n518)));
	assign n547 = (((!i_18_) & (!n833)) + ((i_18_) & (!n833)) + ((i_18_) & (n833)));
	assign n548 = (((!i_19_) & (!n833)) + ((i_19_) & (!n833)) + ((i_19_) & (n833)));
	assign n546 = (((!n93) & (n547) & (!n94) & (n548)) + ((!n93) & (n547) & (n94) & (!n548)) + ((!n93) & (n547) & (n94) & (n548)) + ((n93) & (!n547) & (!n94) & (n548)) + ((n93) & (!n547) & (n94) & (!n548)) + ((n93) & (!n547) & (n94) & (n548)) + ((n93) & (n547) & (!n94) & (n548)) + ((n93) & (n547) & (n94) & (!n548)) + ((n93) & (n547) & (n94) & (n548)));
	assign n550 = (((!i_37_) & (!n970)) + ((!i_37_) & (n970)) + ((i_37_) & (n970)));
	assign n549 = (((!i_30_) & (!i_31_) & (!n550) & (!n688)) + ((!i_30_) & (!i_31_) & (!n550) & (n688)) + ((!i_30_) & (!i_31_) & (n550) & (!n688)) + ((!i_30_) & (!i_31_) & (n550) & (n688)) + ((!i_30_) & (i_31_) & (!n550) & (!n688)) + ((!i_30_) & (i_31_) & (n550) & (!n688)) + ((!i_30_) & (i_31_) & (n550) & (n688)) + ((i_30_) & (!i_31_) & (!n550) & (!n688)) + ((i_30_) & (!i_31_) & (!n550) & (n688)) + ((i_30_) & (!i_31_) & (n550) & (!n688)) + ((i_30_) & (!i_31_) & (n550) & (n688)) + ((i_30_) & (i_31_) & (!n550) & (!n688)) + ((i_30_) & (i_31_) & (!n550) & (n688)) + ((i_30_) & (i_31_) & (n550) & (!n688)) + ((i_30_) & (i_31_) & (n550) & (n688)));
	assign n554 = (((!n371) & (!n522) & (n454)) + ((!n371) & (n522) & (!n454)) + ((!n371) & (n522) & (n454)) + ((n371) & (!n522) & (!n454)) + ((n371) & (!n522) & (n454)) + ((n371) & (n522) & (!n454)) + ((n371) & (n522) & (n454)));
	assign n552 = (((!i_37_) & (!n101) & (!n554)) + ((!i_37_) & (!n101) & (n554)) + ((!i_37_) & (n101) & (!n554)) + ((!i_37_) & (n101) & (n554)) + ((i_37_) & (!n101) & (n554)) + ((i_37_) & (n101) & (!n554)) + ((i_37_) & (n101) & (n554)));
	assign n556 = (((!i_16_) & (n960)) + ((i_16_) & (!n960)) + ((i_16_) & (n960)));
	assign n557 = (((!i_13_) & (!n229)) + ((i_13_) & (!n229)) + ((i_13_) & (n229)));
	assign n558 = (((!i_23_) & (n734)) + ((i_23_) & (!n734)) + ((i_23_) & (n734)));
	assign n559 = (((!i_12_) & (!n229)) + ((i_12_) & (!n229)) + ((i_12_) & (n229)));
	assign n555 = (((!n556) & (n557) & (!n558) & (n559)) + ((!n556) & (n557) & (n558) & (!n559)) + ((!n556) & (n557) & (n558) & (n559)) + ((n556) & (!n557) & (!n558) & (n559)) + ((n556) & (!n557) & (n558) & (!n559)) + ((n556) & (!n557) & (n558) & (n559)) + ((n556) & (n557) & (!n558) & (n559)) + ((n556) & (n557) & (n558) & (!n559)) + ((n556) & (n557) & (n558) & (n559)));
	assign n562 = (((!i_34_) & (!n364) & (!n501) & (!n607)) + ((!i_34_) & (!n364) & (!n501) & (n607)) + ((!i_34_) & (!n364) & (n501) & (!n607)) + ((!i_34_) & (!n364) & (n501) & (n607)) + ((!i_34_) & (n364) & (!n501) & (!n607)) + ((!i_34_) & (n364) & (!n501) & (n607)) + ((!i_34_) & (n364) & (n501) & (!n607)) + ((!i_34_) & (n364) & (n501) & (n607)) + ((i_34_) & (!n364) & (!n501) & (!n607)) + ((i_34_) & (!n364) & (!n501) & (n607)) + ((i_34_) & (!n364) & (n501) & (!n607)) + ((i_34_) & (!n364) & (n501) & (n607)) + ((i_34_) & (n364) & (!n501) & (n607)) + ((i_34_) & (n364) & (n501) & (!n607)) + ((i_34_) & (n364) & (n501) & (n607)));
	assign n561 = (((!i_34_) & (n717)) + ((i_34_) & (!n717)) + ((i_34_) & (n717)));
	assign n560 = (((n562) & (!i_33_) & (!n555) & (n561)) + ((n562) & (!i_33_) & (n555) & (!n561)) + ((n562) & (!i_33_) & (n555) & (n561)) + ((n562) & (i_33_) & (!n555) & (!n561)) + ((n562) & (i_33_) & (!n555) & (n561)) + ((n562) & (i_33_) & (n555) & (!n561)) + ((n562) & (i_33_) & (n555) & (n561)));
	assign n563 = (((n467) & (!n549) & (!n552) & (!n1187)) + ((n467) & (!n549) & (!n552) & (n1187)) + ((n467) & (!n549) & (n552) & (!n1187)) + ((n467) & (!n549) & (n552) & (n1187)) + ((n467) & (n549) & (!n552) & (!n1187)) + ((n467) & (n549) & (!n552) & (n1187)) + ((n467) & (n549) & (n552) & (!n1187)));
	assign n569 = (((n1188) & (!n544) & (!n716) & (n717)) + ((n1188) & (!n544) & (n716) & (!n717)) + ((n1188) & (!n544) & (n716) & (n717)) + ((n1188) & (n544) & (!n716) & (!n717)) + ((n1188) & (n544) & (!n716) & (n717)) + ((n1188) & (n544) & (n716) & (!n717)) + ((n1188) & (n544) & (n716) & (n717)));
	assign n567 = (((!i_30_) & (n560) & (!n563) & (n569)) + ((i_30_) & (!n560) & (!n563) & (n569)) + ((i_30_) & (n560) & (!n563) & (n569)));
	assign n573 = (((!n841) & (!n884)) + ((!n841) & (n884)) + ((n841) & (n884)));
	assign n572 = (((!i_27_) & (!n833)) + ((i_27_) & (!n833)) + ((i_27_) & (n833)));
	assign n570 = (((!n356) & (n573) & (!n572)) + ((!n356) & (n573) & (n572)) + ((n356) & (n573) & (n572)));
	assign n576 = (((!i_8_) & (!n985) & (n586)) + ((!i_8_) & (n985) & (!n586)) + ((!i_8_) & (n985) & (n586)) + ((i_8_) & (!n985) & (!n586)) + ((i_8_) & (!n985) & (n586)) + ((i_8_) & (n985) & (!n586)) + ((i_8_) & (n985) & (n586)));
	assign n575 = (((!i_11_) & (n1010)) + ((i_11_) & (!n1010)) + ((i_11_) & (n1010)));
	assign n574 = (((n576) & (!n70) & (n575)) + ((n576) & (n70) & (!n575)) + ((n576) & (n70) & (n575)));
	assign n578 = (((!n243) & (!n334) & (!i_7_) & (i_28_)) + ((!n243) & (!n334) & (i_7_) & (!i_28_)) + ((!n243) & (!n334) & (i_7_) & (i_28_)) + ((!n243) & (n334) & (!i_7_) & (!i_28_)) + ((!n243) & (n334) & (!i_7_) & (i_28_)) + ((!n243) & (n334) & (i_7_) & (!i_28_)) + ((!n243) & (n334) & (i_7_) & (i_28_)) + ((n243) & (!n334) & (!i_7_) & (!i_28_)) + ((n243) & (!n334) & (!i_7_) & (i_28_)) + ((n243) & (!n334) & (i_7_) & (!i_28_)) + ((n243) & (!n334) & (i_7_) & (i_28_)) + ((n243) & (n334) & (!i_7_) & (!i_28_)) + ((n243) & (n334) & (!i_7_) & (i_28_)) + ((n243) & (n334) & (i_7_) & (!i_28_)) + ((n243) & (n334) & (i_7_) & (i_28_)));
	assign n579 = (((!i_9_) & (!n69) & (!n631) & (!n681) & (!n1016)) + ((!i_9_) & (!n69) & (!n631) & (!n681) & (n1016)) + ((!i_9_) & (!n69) & (!n631) & (n681) & (n1016)) + ((!i_9_) & (!n69) & (n631) & (!n681) & (!n1016)) + ((!i_9_) & (!n69) & (n631) & (!n681) & (n1016)) + ((!i_9_) & (!n69) & (n631) & (n681) & (!n1016)) + ((!i_9_) & (!n69) & (n631) & (n681) & (n1016)) + ((!i_9_) & (n69) & (!n631) & (!n681) & (!n1016)) + ((!i_9_) & (n69) & (!n631) & (!n681) & (n1016)) + ((!i_9_) & (n69) & (!n631) & (n681) & (!n1016)) + ((!i_9_) & (n69) & (!n631) & (n681) & (n1016)) + ((!i_9_) & (n69) & (n631) & (!n681) & (!n1016)) + ((!i_9_) & (n69) & (n631) & (!n681) & (n1016)) + ((!i_9_) & (n69) & (n631) & (n681) & (!n1016)) + ((!i_9_) & (n69) & (n631) & (n681) & (n1016)) + ((i_9_) & (!n69) & (!n631) & (!n681) & (!n1016)) + ((i_9_) & (!n69) & (!n631) & (!n681) & (n1016)) + ((i_9_) & (!n69) & (!n631) & (n681) & (!n1016)) + ((i_9_) & (!n69) & (!n631) & (n681) & (n1016)) + ((i_9_) & (!n69) & (n631) & (!n681) & (!n1016)) + ((i_9_) & (!n69) & (n631) & (!n681) & (n1016)) + ((i_9_) & (!n69) & (n631) & (n681) & (!n1016)) + ((i_9_) & (!n69) & (n631) & (n681) & (n1016)) + ((i_9_) & (n69) & (!n631) & (!n681) & (!n1016)) + ((i_9_) & (n69) & (!n631) & (!n681) & (n1016)) + ((i_9_) & (n69) & (!n631) & (n681) & (!n1016)) + ((i_9_) & (n69) & (!n631) & (n681) & (n1016)) + ((i_9_) & (n69) & (n631) & (!n681) & (!n1016)) + ((i_9_) & (n69) & (n631) & (!n681) & (n1016)) + ((i_9_) & (n69) & (n631) & (n681) & (!n1016)) + ((i_9_) & (n69) & (n631) & (n681) & (n1016)));
	assign n577 = (((n578) & (n579) & (!n570) & (n574)) + ((n578) & (n579) & (n570) & (!n574)) + ((n578) & (n579) & (n570) & (n574)));
	assign n580 = (((!i_10_) & (!i_30_) & (n70) & (!n229)) + ((!i_10_) & (i_30_) & (n70) & (!n229)) + ((!i_10_) & (i_30_) & (n70) & (n229)) + ((i_10_) & (!i_30_) & (!n70) & (!n229)) + ((i_10_) & (!i_30_) & (n70) & (!n229)) + ((i_10_) & (i_30_) & (!n70) & (!n229)) + ((i_10_) & (i_30_) & (!n70) & (n229)) + ((i_10_) & (i_30_) & (n70) & (!n229)) + ((i_10_) & (i_30_) & (n70) & (n229)));
	assign n583 = (((!n442) & (!n580) & (n556)) + ((!n442) & (n580) & (!n556)) + ((!n442) & (n580) & (n556)) + ((n442) & (!n580) & (!n556)) + ((n442) & (!n580) & (n556)) + ((n442) & (n580) & (!n556)) + ((n442) & (n580) & (n556)));
	assign n584 = (((!n543) & (!n973) & (!n993) & (n1186)) + ((!n543) & (!n973) & (n993) & (n1186)) + ((!n543) & (n973) & (!n993) & (n1186)) + ((!n543) & (n973) & (n993) & (n1186)) + ((n543) & (!n973) & (n993) & (n1186)) + ((n543) & (n973) & (!n993) & (n1186)) + ((n543) & (n973) & (n993) & (n1186)));
	assign n582 = (((!i_37_) & (!n577) & (n583) & (n584)) + ((!i_37_) & (n577) & (n583) & (n584)) + ((i_37_) & (n577) & (n583) & (n584)));
	assign n586 = (((!i_18_) & (n1006)) + ((i_18_) & (!n1006)) + ((i_18_) & (n1006)));
	assign n587 = (((!n595) & (n527)) + ((n595) & (!n527)) + ((n595) & (n527)));
	assign n585 = (((!n586) & (!i_8_) & (n587)) + ((!n586) & (i_8_) & (!n587)) + ((!n586) & (i_8_) & (n587)) + ((n586) & (!i_8_) & (!n587)) + ((n586) & (!i_8_) & (n587)) + ((n586) & (i_8_) & (!n587)) + ((n586) & (i_8_) & (n587)));
	assign n590 = (((!i_9_) & (!n575) & (!n585) & (!n1016)) + ((!i_9_) & (!n575) & (!n585) & (n1016)) + ((!i_9_) & (!n575) & (n585) & (!n1016)) + ((!i_9_) & (n575) & (!n585) & (!n1016)) + ((!i_9_) & (n575) & (!n585) & (n1016)));
	assign n588 = (((!i_13_) & (!i_14_) & (!i_33_) & (n590)) + ((!i_13_) & (!i_14_) & (i_33_) & (n590)) + ((!i_13_) & (i_14_) & (!i_33_) & (n590)) + ((i_13_) & (!i_14_) & (!i_33_) & (n590)) + ((i_13_) & (!i_14_) & (i_33_) & (n590)));
	assign n591 = (((!i_33_) & (!n953) & (!n1011) & (!n1016)) + ((!i_33_) & (!n953) & (n1011) & (!n1016)) + ((!i_33_) & (n953) & (!n1011) & (!n1016)) + ((i_33_) & (!n953) & (!n1011) & (!n1016)) + ((i_33_) & (!n953) & (n1011) & (!n1016)));
	assign n595 = (((!i_7_) & (n373)) + ((i_7_) & (!n373)) + ((i_7_) & (n373)));
	assign n594 = (((!n522) & (!n595) & (n550)) + ((!n522) & (n595) & (!n550)) + ((!n522) & (n595) & (n550)) + ((n522) & (!n595) & (!n550)) + ((n522) & (!n595) & (n550)) + ((n522) & (n595) & (!n550)) + ((n522) & (n595) & (n550)));
	assign n596 = (((!n521) & (!n594) & (!n622) & (!n965)) + ((!n521) & (!n594) & (!n622) & (n965)) + ((!n521) & (n594) & (!n622) & (!n965)) + ((n521) & (!n594) & (!n622) & (!n965)) + ((n521) & (!n594) & (!n622) & (n965)));
	assign n601 = (((!i_37_) & (!n588) & (!n591) & (!n596)) + ((!i_37_) & (!n588) & (n591) & (!n596)) + ((!i_37_) & (n588) & (!n591) & (!n596)) + ((!i_37_) & (n588) & (n591) & (!n596)) + ((i_37_) & (!n588) & (!n591) & (!n596)));
	assign n607 = (((!i_8_) & (!n15)) + ((i_8_) & (!n15)) + ((i_8_) & (n15)));
	assign n608 = (((!i_17_) & (!n833)) + ((i_17_) & (!n833)) + ((i_17_) & (n833)));
	assign n609 = (((!i_8_) & (n734)) + ((i_8_) & (!n734)) + ((i_8_) & (n734)));
	assign n605 = (((!n364) & (!n607) & (!n608) & (n609)) + ((!n364) & (!n607) & (n608) & (!n609)) + ((!n364) & (!n607) & (n608) & (n609)) + ((!n364) & (n607) & (!n608) & (n609)) + ((!n364) & (n607) & (n608) & (!n609)) + ((!n364) & (n607) & (n608) & (n609)) + ((n364) & (n607) & (!n608) & (n609)) + ((n364) & (n607) & (n608) & (!n609)) + ((n364) & (n607) & (n608) & (n609)));
	assign n611 = (((!i_33_) & (n974)) + ((i_33_) & (!n974)) + ((i_33_) & (n974)));
	assign n612 = (((n789) & (n1259)));
	assign n610 = (((!n605) & (n611) & (!n612) & (n241)) + ((!n605) & (n611) & (n612) & (!n241)) + ((!n605) & (n611) & (n612) & (n241)) + ((n605) & (!n611) & (!n612) & (n241)) + ((n605) & (!n611) & (n612) & (!n241)) + ((n605) & (!n611) & (n612) & (n241)) + ((n605) & (n611) & (!n612) & (n241)) + ((n605) & (n611) & (n612) & (!n241)) + ((n605) & (n611) & (n612) & (n241)));
	assign n614 = (((!n689) & (!n953)) + ((!n689) & (n953)) + ((n689) & (n953)));
	assign n615 = (((!i_29_) & (!n601) & (!n1027) & (n1256)) + ((!i_29_) & (!n601) & (n1027) & (n1256)) + ((!i_29_) & (n601) & (!n1027) & (n1256)) + ((!i_29_) & (n601) & (n1027) & (n1256)) + ((i_29_) & (!n601) & (n1027) & (n1256)) + ((i_29_) & (n601) & (!n1027) & (n1256)) + ((i_29_) & (n601) & (n1027) & (n1256)));
	assign n613 = (((!n543) & (!n610) & (n614) & (n615)) + ((!n543) & (n610) & (n614) & (n615)) + ((n543) & (n610) & (n614) & (n615)));
	assign n617 = (((!i_25_) & (!i_28_) & (!n497) & (!n1026)) + ((!i_25_) & (!i_28_) & (!n497) & (n1026)) + ((!i_25_) & (!i_28_) & (n497) & (!n1026)) + ((!i_25_) & (!i_28_) & (n497) & (n1026)) + ((!i_25_) & (i_28_) & (!n497) & (!n1026)) + ((!i_25_) & (i_28_) & (!n497) & (n1026)) + ((!i_25_) & (i_28_) & (n497) & (!n1026)) + ((!i_25_) & (i_28_) & (n497) & (n1026)) + ((i_25_) & (!i_28_) & (!n497) & (n1026)) + ((i_25_) & (!i_28_) & (n497) & (!n1026)) + ((i_25_) & (!i_28_) & (n497) & (n1026)) + ((i_25_) & (i_28_) & (!n497) & (!n1026)) + ((i_25_) & (i_28_) & (!n497) & (n1026)) + ((i_25_) & (i_28_) & (n497) & (!n1026)) + ((i_25_) & (i_28_) & (n497) & (n1026)));
	assign n616 = (((!n404) & (!n501) & (!n609) & (n617)) + ((!n404) & (!n501) & (n609) & (n617)) + ((!n404) & (n501) & (!n609) & (n617)) + ((!n404) & (n501) & (n609) & (n617)) + ((n404) & (!n501) & (n609) & (n617)) + ((n404) & (n501) & (!n609) & (n617)) + ((n404) & (n501) & (n609) & (n617)));
	assign n619 = (((!i_8_) & (n1030)) + ((i_8_) & (!n1030)) + ((i_8_) & (n1030)));
	assign n620 = (((!i_8_) & (n735)) + ((i_8_) & (!n735)) + ((i_8_) & (n735)));
	assign n618 = (((!n364) & (!n608) & (!n619) & (n620)) + ((!n364) & (!n608) & (n619) & (n620)) + ((!n364) & (n608) & (!n619) & (!n620)) + ((!n364) & (n608) & (!n619) & (n620)) + ((!n364) & (n608) & (n619) & (!n620)) + ((!n364) & (n608) & (n619) & (n620)) + ((n364) & (!n608) & (n619) & (n620)) + ((n364) & (n608) & (n619) & (!n620)) + ((n364) & (n608) & (n619) & (n620)));
	assign n623 = (((!i_10_) & (!n1016) & (!i_33_) & (i_9_)) + ((!i_10_) & (!n1016) & (i_33_) & (!i_9_)) + ((!i_10_) & (!n1016) & (i_33_) & (i_9_)) + ((!i_10_) & (n1016) & (!i_33_) & (!i_9_)) + ((!i_10_) & (n1016) & (!i_33_) & (i_9_)) + ((!i_10_) & (n1016) & (i_33_) & (!i_9_)) + ((!i_10_) & (n1016) & (i_33_) & (i_9_)) + ((i_10_) & (!n1016) & (!i_33_) & (!i_9_)) + ((i_10_) & (!n1016) & (!i_33_) & (i_9_)) + ((i_10_) & (!n1016) & (i_33_) & (!i_9_)) + ((i_10_) & (!n1016) & (i_33_) & (i_9_)) + ((i_10_) & (n1016) & (!i_33_) & (!i_9_)) + ((i_10_) & (n1016) & (!i_33_) & (i_9_)) + ((i_10_) & (n1016) & (i_33_) & (!i_9_)) + ((i_10_) & (n1016) & (i_33_) & (i_9_)));
	assign n622 = (((!i_1_) & (n1007)) + ((i_1_) & (!n1007)) + ((i_1_) & (n1007)));
	assign n621 = (((n623) & (!n373) & (!n101) & (n622)) + ((n623) & (!n373) & (n101) & (!n622)) + ((n623) & (!n373) & (n101) & (n622)) + ((n623) & (n373) & (!n101) & (!n622)) + ((n623) & (n373) & (!n101) & (n622)) + ((n623) & (n373) & (n101) & (!n622)) + ((n623) & (n373) & (n101) & (n622)));
	assign n626 = (((!n461) & (!n467) & (!n550)) + ((!n461) & (!n467) & (n550)) + ((!n461) & (n467) & (n550)) + ((n461) & (!n467) & (!n550)) + ((n461) & (!n467) & (n550)) + ((n461) & (n467) & (!n550)) + ((n461) & (n467) & (n550)));
	assign n624 = (((!i_37_) & (!n621) & (n626) & (!n681)) + ((!i_37_) & (!n621) & (n626) & (n681)) + ((!i_37_) & (n621) & (n626) & (!n681)) + ((!i_37_) & (n621) & (n626) & (n681)) + ((i_37_) & (!n621) & (n626) & (!n681)) + ((i_37_) & (n621) & (n626) & (!n681)) + ((i_37_) & (n621) & (n626) & (n681)));
	assign n628 = (((!i_20_) & (n734)) + ((i_20_) & (!n734)) + ((i_20_) & (n734)));
	assign n629 = (((!i_20_) & (n735)) + ((i_20_) & (!n735)) + ((i_20_) & (n735)));
	assign n627 = (((!n501) & (!n543) & (n628) & (!n629)) + ((!n501) & (!n543) & (n628) & (n629)) + ((!n501) & (n543) & (n628) & (n629)) + ((n501) & (!n543) & (!n628) & (!n629)) + ((n501) & (!n543) & (!n628) & (n629)) + ((n501) & (!n543) & (n628) & (!n629)) + ((n501) & (!n543) & (n628) & (n629)) + ((n501) & (n543) & (!n628) & (n629)) + ((n501) & (n543) & (n628) & (n629)));
	assign n631 = (((!i_20_) & (n1006)) + ((i_20_) & (!n1006)) + ((i_20_) & (n1006)));
	assign n630 = (((!i_12_) & (n627) & (!n500) & (n631)) + ((!i_12_) & (n627) & (n500) & (!n631)) + ((!i_12_) & (n627) & (n500) & (n631)) + ((i_12_) & (!n627) & (!n500) & (n631)) + ((i_12_) & (!n627) & (n500) & (!n631)) + ((i_12_) & (!n627) & (n500) & (n631)) + ((i_12_) & (n627) & (!n500) & (n631)) + ((i_12_) & (n627) & (n500) & (!n631)) + ((i_12_) & (n627) & (n500) & (n631)));
	assign n632 = (((!i_7_) & (i_37_) & (n349)));
	assign n633 = (((n350) & (!n632) & (i_25_) & (n246)) + ((n350) & (n632) & (!i_25_) & (!n246)) + ((n350) & (n632) & (!i_25_) & (n246)) + ((n350) & (n632) & (i_25_) & (!n246)) + ((n350) & (n632) & (i_25_) & (n246)));
	assign n634 = (((!n253) & (!n531) & (!n633) & (!n954)) + ((!n253) & (!n531) & (!n633) & (n954)) + ((!n253) & (n531) & (!n633) & (!n954)) + ((!n253) & (n531) & (!n633) & (n954)) + ((n253) & (!n531) & (!n633) & (!n954)) + ((n253) & (!n531) & (!n633) & (n954)) + ((n253) & (n531) & (!n633) & (!n954)));
	assign n639 = (((!i_9_) & (n735)) + ((i_9_) & (!n735)) + ((i_9_) & (n735)));
	assign n640 = (((!i_9_) & (n734)) + ((i_9_) & (!n734)) + ((i_9_) & (n734)));
	assign n638 = (((!n501) & (!n543) & (!n639) & (n640)) + ((!n501) & (!n543) & (n639) & (n640)) + ((!n501) & (n543) & (n639) & (n640)) + ((n501) & (!n543) & (!n639) & (!n640)) + ((n501) & (!n543) & (!n639) & (n640)) + ((n501) & (!n543) & (n639) & (!n640)) + ((n501) & (!n543) & (n639) & (n640)) + ((n501) & (n543) & (n639) & (!n640)) + ((n501) & (n543) & (n639) & (n640)));
	assign n641 = (((!n544) & (n443) & (!n448) & (n534)) + ((!n544) & (n443) & (n448) & (!n534)) + ((!n544) & (n443) & (n448) & (n534)) + ((n544) & (!n443) & (!n448) & (n534)) + ((n544) & (!n443) & (n448) & (!n534)) + ((n544) & (!n443) & (n448) & (n534)) + ((n544) & (n443) & (!n448) & (n534)) + ((n544) & (n443) & (n448) & (!n534)) + ((n544) & (n443) & (n448) & (n534)));
	assign n644 = (((!n986) & (n1011)) + ((n986) & (!n1011)) + ((n986) & (n1011)));
	assign n643 = (((!i_11_) & (!n70) & (n1010)) + ((!i_11_) & (n70) & (!n1010)) + ((!i_11_) & (n70) & (n1010)) + ((i_11_) & (!n70) & (!n1010)) + ((i_11_) & (!n70) & (n1010)) + ((i_11_) & (n70) & (!n1010)) + ((i_11_) & (n70) & (n1010)));
	assign n642 = (((n644) & (!i_13_) & (n643) & (n576)) + ((n644) & (i_13_) & (!n643) & (!n576)) + ((n644) & (i_13_) & (!n643) & (n576)) + ((n644) & (i_13_) & (n643) & (!n576)) + ((n644) & (i_13_) & (n643) & (n576)));
	assign n646 = (((!n63) & (n522)) + ((n63) & (!n522)) + ((n63) & (n522)));
	assign n645 = (((!n642) & (n443) & (!n448) & (n646)) + ((!n642) & (n443) & (n448) & (!n646)) + ((!n642) & (n443) & (n448) & (n646)) + ((n642) & (!n443) & (!n448) & (n646)) + ((n642) & (!n443) & (n448) & (!n646)) + ((n642) & (!n443) & (n448) & (n646)) + ((n642) & (n443) & (!n448) & (n646)) + ((n642) & (n443) & (n448) & (!n646)) + ((n642) & (n443) & (n448) & (n646)));
	assign n648 = (((!i_32_) & (n978)) + ((i_32_) & (!n978)) + ((i_32_) & (n978)));
	assign n649 = (((!i_24_) & (n1004)) + ((i_24_) & (!n1004)) + ((i_24_) & (n1004)));
	assign n647 = (((!n334) & (!n362) & (!n648) & (n649)) + ((!n334) & (!n362) & (n648) & (!n649)) + ((!n334) & (!n362) & (n648) & (n649)) + ((n334) & (!n362) & (!n648) & (n649)) + ((n334) & (!n362) & (n648) & (!n649)) + ((n334) & (!n362) & (n648) & (n649)) + ((n334) & (n362) & (!n648) & (n649)) + ((n334) & (n362) & (n648) & (!n649)) + ((n334) & (n362) & (n648) & (n649)));
	assign n651 = (((n1179) & (!n984) & (!n639) & (n1013)) + ((n1179) & (!n984) & (n639) & (!n1013)) + ((n1179) & (!n984) & (n639) & (n1013)) + ((n1179) & (n984) & (!n639) & (!n1013)) + ((n1179) & (n984) & (!n639) & (n1013)) + ((n1179) & (n984) & (n639) & (!n1013)) + ((n1179) & (n984) & (n639) & (n1013)));
	assign n650 = (((n651) & (!n66) & (!n515) & (n469)) + ((n651) & (!n66) & (n515) & (!n469)) + ((n651) & (!n66) & (n515) & (n469)) + ((n651) & (n66) & (!n515) & (!n469)) + ((n651) & (n66) & (!n515) & (n469)) + ((n651) & (n66) & (n515) & (!n469)) + ((n651) & (n66) & (n515) & (n469)));
	assign n653 = (((!n367) & (!n572)) + ((!n367) & (n572)) + ((n367) & (n572)));
	assign n654 = (((!n59) & (n505)) + ((n59) & (!n505)) + ((n59) & (n505)));
	assign n652 = (((!n404) & (!n554) & (n653) & (!n654)) + ((!n404) & (!n554) & (n653) & (n654)) + ((!n404) & (n554) & (!n653) & (!n654)) + ((!n404) & (n554) & (!n653) & (n654)) + ((!n404) & (n554) & (n653) & (!n654)) + ((!n404) & (n554) & (n653) & (n654)) + ((n404) & (!n554) & (n653) & (n654)) + ((n404) & (n554) & (!n653) & (n654)) + ((n404) & (n554) & (n653) & (n654)));
	assign n657 = (((!n215) & (!n367)) + ((n215) & (!n367)) + ((n215) & (n367)));
	assign n655 = (((!n349) & (!n376) & (!n404) & (!n657)) + ((!n349) & (!n376) & (!n404) & (n657)) + ((!n349) & (n376) & (!n404) & (!n657)) + ((!n349) & (n376) & (!n404) & (n657)) + ((!n349) & (n376) & (n404) & (!n657)) + ((!n349) & (n376) & (n404) & (n657)) + ((n349) & (!n376) & (!n404) & (n657)) + ((n349) & (n376) & (!n404) & (n657)) + ((n349) & (n376) & (n404) & (n657)));
	assign n660 = (((!n652) & (n988) & (!n647) & (n650)) + ((!n652) & (n988) & (n647) & (!n650)) + ((!n652) & (n988) & (n647) & (n650)) + ((n652) & (!n988) & (!n647) & (n650)) + ((n652) & (!n988) & (n647) & (!n650)) + ((n652) & (!n988) & (n647) & (n650)) + ((n652) & (n988) & (!n647) & (n650)) + ((n652) & (n988) & (n647) & (!n650)) + ((n652) & (n988) & (n647) & (n650)));
	assign n661 = (((n1180) & (n1181) & (!n655) & (n1029)) + ((n1180) & (n1181) & (n655) & (!n1029)) + ((n1180) & (n1181) & (n655) & (n1029)));
	assign n659 = (((!n986) & (n953)) + ((n986) & (!n953)) + ((n986) & (n953)));
	assign n658 = (((n660) & (n661) & (!n570) & (n659)) + ((n660) & (n661) & (n570) & (!n659)) + ((n660) & (n661) & (n570) & (n659)));
	assign n664 = (((!i_26_) & (n1004)) + ((i_26_) & (!n1004)) + ((i_26_) & (n1004)));
	assign n662 = (((!i_33_) & (!n245) & (!n362) & (!n664)) + ((!i_33_) & (!n245) & (!n362) & (n664)) + ((!i_33_) & (!n245) & (n362) & (!n664)) + ((!i_33_) & (!n245) & (n362) & (n664)) + ((!i_33_) & (n245) & (!n362) & (!n664)) + ((!i_33_) & (n245) & (!n362) & (n664)) + ((i_33_) & (!n245) & (!n362) & (n664)) + ((i_33_) & (!n245) & (n362) & (n664)) + ((i_33_) & (n245) & (!n362) & (n664)));
	assign n665 = (((i_20_) & (!i_23_) & (i_25_) & (!n849)));
	assign n670 = (((!i_34_) & (n531)));
	assign n668 = (((!i_27_) & (n891)));
	assign n669 = (((i_22_) & (n1024)));
	assign n667 = (((i_35_) & (n670) & (!n668) & (n669)) + ((i_35_) & (n670) & (n668) & (!n669)) + ((i_35_) & (n670) & (n668) & (n669)));
	assign n672 = (((i_25_) & (n1024)));
	assign n673 = (((n350) & (i_33_)));
	assign n671 = (((n253) & (!n665) & (n672) & (n673)) + ((n253) & (n665) & (!n672) & (!n673)) + ((n253) & (n665) & (!n672) & (n673)) + ((n253) & (n665) & (n672) & (!n673)) + ((n253) & (n665) & (n672) & (n673)));
	assign n676 = (((!i_34_) & (!n494) & (!n880) & (n1175)) + ((!i_34_) & (!n494) & (n880) & (n1175)) + ((!i_34_) & (n494) & (!n880) & (n1175)) + ((!i_34_) & (n494) & (n880) & (n1175)) + ((i_34_) & (!n494) & (!n880) & (n1175)) + ((i_34_) & (!n494) & (n880) & (n1175)) + ((i_34_) & (n494) & (!n880) & (n1175)));
	assign n674 = (((!n498) & (n662) & (!n671) & (n676)) + ((n498) & (!n662) & (!n671) & (n676)) + ((n498) & (n662) & (!n671) & (n676)));
	assign n677 = (((i_34_) & (n494) & (!n522)));
	assign n680 = (((!i_20_) & (!i_21_)));
	assign n681 = (((n467) & (n494)));
	assign n682 = (((!n953) & (!n1011)) + ((!n953) & (n1011)) + ((n953) & (!n1011)));
	assign n679 = (((n680) & (i_2_) & (n681) & (n682)));
	assign n684 = (((!i_34_) & (n163)) + ((i_34_) & (!n163)) + ((i_34_) & (n163)));
	assign n685 = (((!i_31_) & (i_32_)) + ((i_31_) & (!i_32_)) + ((i_31_) & (i_32_)));
	assign n683 = (((!i_22_) & (!n684) & (!n685) & (!n692)) + ((!i_22_) & (!n684) & (!n685) & (n692)) + ((!i_22_) & (!n684) & (n685) & (!n692)) + ((!i_22_) & (!n684) & (n685) & (n692)) + ((!i_22_) & (n684) & (!n685) & (!n692)) + ((!i_22_) & (n684) & (!n685) & (n692)) + ((!i_22_) & (n684) & (n685) & (!n692)) + ((!i_22_) & (n684) & (n685) & (n692)) + ((i_22_) & (!n684) & (!n685) & (!n692)) + ((i_22_) & (!n684) & (n685) & (!n692)) + ((i_22_) & (!n684) & (n685) & (n692)) + ((i_22_) & (n684) & (!n685) & (!n692)) + ((i_22_) & (n684) & (!n685) & (n692)) + ((i_22_) & (n684) & (n685) & (!n692)) + ((i_22_) & (n684) & (n685) & (n692)));
	assign n689 = (((i_29_) & (n495)));
	assign n688 = (((!n522) & (!n1011)) + ((!n522) & (n1011)) + ((n522) & (!n1011)));
	assign n686 = (((!n453) & (!n664) & (n689) & (!n688)) + ((!n453) & (!n664) & (n689) & (n688)) + ((n453) & (!n664) & (n689) & (n688)));
	assign n692 = (((!i_30_) & (n531)));
	assign n691 = (((n495) & (!n677) & (n692) & (!n973)) + ((n495) & (n677) & (!n692) & (!n973)) + ((n495) & (n677) & (!n692) & (n973)) + ((n495) & (n677) & (n692) & (!n973)) + ((n495) & (n677) & (n692) & (n973)));
	assign n695 = (((!n96) & (n522)) + ((n96) & (!n522)) + ((n96) & (n522)));
	assign n696 = (((!n96) & (n609)) + ((n96) & (!n609)) + ((n96) & (n609)));
	assign n694 = (((!n404) & (!n653) & (n695) & (!n696)) + ((!n404) & (!n653) & (n695) & (n696)) + ((!n404) & (n653) & (!n695) & (!n696)) + ((!n404) & (n653) & (!n695) & (n696)) + ((!n404) & (n653) & (n695) & (!n696)) + ((!n404) & (n653) & (n695) & (n696)) + ((n404) & (!n653) & (n695) & (n696)) + ((n404) & (n653) & (!n695) & (n696)) + ((n404) & (n653) & (n695) & (n696)));
	assign n698 = (((n1174) & (!n555) & (!n611) & (n649)) + ((n1174) & (!n555) & (n611) & (!n649)) + ((n1174) & (!n555) & (n611) & (n649)) + ((n1174) & (n555) & (!n611) & (!n649)) + ((n1174) & (n555) & (!n611) & (n649)) + ((n1174) & (n555) & (n611) & (!n649)) + ((n1174) & (n555) & (n611) & (n649)));
	assign n699 = (((!n404) & (!n653) & (!n1021) & (n1023)) + ((!n404) & (!n653) & (n1021) & (n1023)) + ((!n404) & (n653) & (!n1021) & (!n1023)) + ((!n404) & (n653) & (!n1021) & (n1023)) + ((!n404) & (n653) & (n1021) & (!n1023)) + ((!n404) & (n653) & (n1021) & (n1023)) + ((n404) & (!n653) & (n1021) & (n1023)) + ((n404) & (n653) & (n1021) & (!n1023)) + ((n404) & (n653) & (n1021) & (n1023)));
	assign n697 = (((n698) & (n699) & (!i_33_) & (n694)) + ((n698) & (n699) & (i_33_) & (!n694)) + ((n698) & (n699) & (i_33_) & (n694)));
	assign n700 = (((!i_28_) & (!n376) & (!n833)) + ((!i_28_) & (n376) & (!n833)) + ((!i_28_) & (n376) & (n833)) + ((i_28_) & (!n376) & (!n833)) + ((i_28_) & (!n376) & (n833)) + ((i_28_) & (n376) & (!n833)) + ((i_28_) & (n376) & (n833)));
	assign n703 = (((n1260) & (n517)));
	assign n704 = (((!i_14_) & (!n1014) & (n556)) + ((!i_14_) & (n1014) & (!n556)) + ((!i_14_) & (n1014) & (n556)) + ((i_14_) & (!n1014) & (!n556)) + ((i_14_) & (!n1014) & (n556)) + ((i_14_) & (n1014) & (!n556)) + ((i_14_) & (n1014) & (n556)));
	assign n702 = (((!n703) & (n345) & (!n648) & (n704)) + ((!n703) & (n345) & (n648) & (!n704)) + ((!n703) & (n345) & (n648) & (n704)) + ((n703) & (!n345) & (!n648) & (n704)) + ((n703) & (!n345) & (n648) & (!n704)) + ((n703) & (!n345) & (n648) & (n704)) + ((n703) & (n345) & (!n648) & (n704)) + ((n703) & (n345) & (n648) & (!n704)) + ((n703) & (n345) & (n648) & (n704)));
	assign n705 = (((!n121) & (!n243) & (!n700) & (!n716)) + ((!n121) & (!n243) & (!n700) & (n716)) + ((n121) & (!n243) & (!n700) & (!n716)) + ((n121) & (!n243) & (!n700) & (n716)) + ((n121) & (!n243) & (n700) & (!n716)));
	assign n710 = (((!n356) & (!n572) & (!n1022)) + ((!n356) & (!n572) & (n1022)) + ((!n356) & (n572) & (!n1022)) + ((!n356) & (n572) & (n1022)) + ((n356) & (!n572) & (n1022)) + ((n356) & (n572) & (!n1022)) + ((n356) & (n572) & (n1022)));
	assign n709 = (((!n649) & (n702) & (!n705) & (n710)) + ((n649) & (!n702) & (!n705) & (n710)) + ((n649) & (n702) & (!n705) & (n710)));
	assign n712 = (((!n347) & (!n367) & (!n480) & (n696)) + ((!n347) & (!n367) & (n480) & (n696)) + ((!n347) & (n367) & (n480) & (n696)) + ((n347) & (!n367) & (!n480) & (!n696)) + ((n347) & (!n367) & (!n480) & (n696)) + ((n347) & (!n367) & (n480) & (!n696)) + ((n347) & (!n367) & (n480) & (n696)) + ((n347) & (n367) & (n480) & (!n696)) + ((n347) & (n367) & (n480) & (n696)));
	assign n714 = (((!n350) & (!n561) & (!n1021)) + ((!n350) & (!n561) & (n1021)) + ((!n350) & (n561) & (!n1021)) + ((!n350) & (n561) & (n1021)) + ((n350) & (!n561) & (n1021)) + ((n350) & (n561) & (!n1021)) + ((n350) & (n561) & (n1021)));
	assign n713 = (((n714) & (!n712) & (n446)) + ((n714) & (n712) & (!n446)) + ((n714) & (n712) & (n446)));
	assign n718 = (((!i_37_) & (!n334) & (!n479)) + ((!i_37_) & (!n334) & (n479)) + ((!i_37_) & (n334) & (!n479)) + ((!i_37_) & (n334) & (n479)) + ((i_37_) & (!n334) & (n479)) + ((i_37_) & (n334) & (!n479)) + ((i_37_) & (n334) & (n479)));
	assign n716 = (((!i_34_) & (n970)) + ((i_34_) & (!n970)) + ((i_34_) & (n970)));
	assign n717 = (((!i_35_) & (!i_37_)) + ((!i_35_) & (i_37_)) + ((i_35_) & (!i_37_)));
	assign n715 = (((!n688) & (n718) & (!n716) & (!n717)) + ((!n688) & (n718) & (!n716) & (n717)) + ((!n688) & (n718) & (n716) & (!n717)) + ((!n688) & (n718) & (n716) & (n717)) + ((n688) & (n718) & (!n716) & (n717)) + ((n688) & (n718) & (n716) & (!n717)) + ((n688) & (n718) & (n716) & (n717)));
	assign n720 = (((!n460) & (!n467) & (!n628)) + ((!n460) & (!n467) & (n628)) + ((!n460) & (n467) & (n628)) + ((n460) & (!n467) & (!n628)) + ((n460) & (!n467) & (n628)) + ((n460) & (n467) & (!n628)) + ((n460) & (n467) & (n628)));
	assign n721 = (((!n640) & (!n1009) & (n587)) + ((!n640) & (n1009) & (!n587)) + ((!n640) & (n1009) & (n587)) + ((n640) & (!n1009) & (!n587)) + ((n640) & (!n1009) & (n587)) + ((n640) & (n1009) & (!n587)) + ((n640) & (n1009) & (n587)));
	assign n719 = (((n720) & (n721) & (!n518) & (n470)) + ((n720) & (n721) & (n518) & (!n470)) + ((n720) & (n721) & (n518) & (n470)));
	assign n723 = (((!i_27_) & (n995)) + ((i_27_) & (!n995)) + ((i_27_) & (n995)));
	assign n724 = (((!i_31_) & (!i_34_)) + ((!i_31_) & (i_34_)) + ((i_31_) & (!i_34_)));
	assign n722 = (((!n253) & (!n649) & (!n723) & (n724)) + ((!n253) & (!n649) & (n723) & (n724)) + ((!n253) & (n649) & (!n723) & (!n724)) + ((!n253) & (n649) & (!n723) & (n724)) + ((!n253) & (n649) & (n723) & (!n724)) + ((!n253) & (n649) & (n723) & (n724)) + ((n253) & (!n649) & (n723) & (n724)) + ((n253) & (n649) & (n723) & (!n724)) + ((n253) & (n649) & (n723) & (n724)));
	assign n725 = (((!i_31_) & (!n362) & (!n664) & (!n724)) + ((!i_31_) & (!n362) & (!n664) & (n724)) + ((!i_31_) & (!n362) & (n664) & (!n724)) + ((!i_31_) & (!n362) & (n664) & (n724)) + ((!i_31_) & (n362) & (!n664) & (n724)) + ((!i_31_) & (n362) & (n664) & (n724)) + ((i_31_) & (!n362) & (n664) & (!n724)) + ((i_31_) & (!n362) & (n664) & (n724)) + ((i_31_) & (n362) & (n664) & (n724)));
	assign n727 = (((!n215) & (!n253) & (!n315)) + ((!n215) & (!n253) & (n315)) + ((!n215) & (n253) & (n315)) + ((n215) & (!n253) & (!n315)) + ((n215) & (!n253) & (n315)) + ((n215) & (n253) & (!n315)) + ((n215) & (n253) & (n315)));
	assign n728 = (((!i_20_) & (!n722) & (!n960)) + ((!i_20_) & (!n722) & (n960)) + ((!i_20_) & (n722) & (!n960)) + ((!i_20_) & (n722) & (n960)) + ((i_20_) & (!n722) & (n960)) + ((i_20_) & (n722) & (!n960)) + ((i_20_) & (n722) & (n960)));
	assign n726 = (((n727) & (n728) & (!n725) & (n608)) + ((n727) & (n728) & (n725) & (!n608)) + ((n727) & (n728) & (n725) & (n608)));
	assign n729 = (((n364) & (!n725)));
	assign n731 = (((!n15) & (!n729) & (!n1030) & (!n1170)) + ((!n15) & (n729) & (!n1030) & (!n1170)) + ((!n15) & (n729) & (!n1030) & (n1170)) + ((n15) & (!n729) & (!n1030) & (!n1170)) + ((n15) & (!n729) & (n1030) & (!n1170)) + ((n15) & (n729) & (!n1030) & (!n1170)) + ((n15) & (n729) & (!n1030) & (n1170)) + ((n15) & (n729) & (n1030) & (!n1170)) + ((n15) & (n729) & (n1030) & (n1170)));
	assign n734 = (((!i_16_) & (i_13_)) + ((i_16_) & (!i_13_)) + ((i_16_) & (i_13_)));
	assign n735 = (((!i_16_) & (i_14_)) + ((i_16_) & (!i_14_)) + ((i_16_) & (i_14_)));
	assign n733 = (((!n726) & (!n731) & (n734) & (n735)) + ((n726) & (!n731) & (!n734) & (!n735)) + ((n726) & (!n731) & (!n734) & (n735)) + ((n726) & (!n731) & (n734) & (!n735)) + ((n726) & (!n731) & (n734) & (n735)));
	assign n739 = (((!n138) & (!n497) & (!i_34_) & (i_24_)) + ((!n138) & (!n497) & (i_34_) & (!i_24_)) + ((!n138) & (!n497) & (i_34_) & (i_24_)) + ((!n138) & (n497) & (!i_34_) & (!i_24_)) + ((!n138) & (n497) & (!i_34_) & (i_24_)) + ((!n138) & (n497) & (i_34_) & (!i_24_)) + ((!n138) & (n497) & (i_34_) & (i_24_)) + ((n138) & (!n497) & (!i_34_) & (!i_24_)) + ((n138) & (!n497) & (!i_34_) & (i_24_)) + ((n138) & (!n497) & (i_34_) & (!i_24_)) + ((n138) & (!n497) & (i_34_) & (i_24_)) + ((n138) & (n497) & (!i_34_) & (!i_24_)) + ((n138) & (n497) & (!i_34_) & (i_24_)) + ((n138) & (n497) & (i_34_) & (!i_24_)) + ((n138) & (n497) & (i_34_) & (i_24_)));
	assign n737 = (((!i_28_) & (!n246) & (!n290) & (n739)) + ((!i_28_) & (!n246) & (n290) & (n739)) + ((!i_28_) & (n246) & (!n290) & (n739)) + ((i_28_) & (!n246) & (!n290) & (n739)) + ((i_28_) & (!n246) & (n290) & (n739)) + ((i_28_) & (n246) & (!n290) & (n739)) + ((i_28_) & (n246) & (n290) & (n739)));
	assign n741 = (((!n11) & (!n684)) + ((!n11) & (n684)) + ((n11) & (n684)));
	assign n740 = (((!i_20_) & (!n497) & (!n737) & (n741)) + ((!i_20_) & (!n497) & (n737) & (n741)) + ((!i_20_) & (n497) & (!n737) & (!n741)) + ((!i_20_) & (n497) & (!n737) & (n741)) + ((!i_20_) & (n497) & (n737) & (!n741)) + ((!i_20_) & (n497) & (n737) & (n741)) + ((i_20_) & (!n497) & (n737) & (n741)) + ((i_20_) & (n497) & (n737) & (!n741)) + ((i_20_) & (n497) & (n737) & (n741)));
	assign n743 = (((!n514) & (n444) & (!n452) & (n653)) + ((!n514) & (n444) & (n452) & (!n653)) + ((!n514) & (n444) & (n452) & (n653)) + ((n514) & (!n444) & (!n452) & (n653)) + ((n514) & (!n444) & (n452) & (!n653)) + ((n514) & (!n444) & (n452) & (n653)) + ((n514) & (n444) & (!n452) & (n653)) + ((n514) & (n444) & (n452) & (!n653)) + ((n514) & (n444) & (n452) & (n653)));
	assign n744 = (((!n469) & (!n501) & (n518) & (!n543)) + ((!n469) & (n501) & (!n518) & (!n543)) + ((!n469) & (n501) & (n518) & (!n543)) + ((n469) & (!n501) & (n518) & (!n543)) + ((n469) & (!n501) & (n518) & (n543)) + ((n469) & (n501) & (!n518) & (!n543)) + ((n469) & (n501) & (!n518) & (n543)) + ((n469) & (n501) & (n518) & (!n543)) + ((n469) & (n501) & (n518) & (n543)));
	assign n747 = (((!n627) & (!n681) & (!n975)) + ((!n627) & (!n681) & (n975)) + ((!n627) & (n681) & (n975)) + ((n627) & (!n681) & (!n975)) + ((n627) & (!n681) & (n975)) + ((n627) & (n681) & (!n975)) + ((n627) & (n681) & (n975)));
	assign n746 = (((!i_19_) & (n1008)) + ((i_19_) & (!n1008)) + ((i_19_) & (n1008)));
	assign n745 = (((n747) & (!n744) & (!n84) & (n746)) + ((n747) & (!n744) & (n84) & (!n746)) + ((n747) & (!n744) & (n84) & (n746)) + ((n747) & (n744) & (!n84) & (!n746)) + ((n747) & (n744) & (!n84) & (n746)) + ((n747) & (n744) & (n84) & (!n746)) + ((n747) & (n744) & (n84) & (n746)));
	assign n749 = (((!i_14_) & (!n40) & (!n364)) + ((!i_14_) & (n40) & (!n364)) + ((!i_14_) & (n40) & (n364)) + ((i_14_) & (!n40) & (!n364)) + ((i_14_) & (!n40) & (n364)) + ((i_14_) & (n40) & (!n364)) + ((i_14_) & (n40) & (n364)));
	assign n748 = (((n749) & (!n546) & (n453)) + ((n749) & (n546) & (!n453)) + ((n749) & (n546) & (n453)));
	assign n750 = (((!i_30_) & (!i_34_) & (!n616) & (!n1182)) + ((!i_30_) & (!i_34_) & (n616) & (!n1182)) + ((!i_30_) & (i_34_) & (!n616) & (!n1182)) + ((!i_30_) & (i_34_) & (!n616) & (n1182)) + ((!i_30_) & (i_34_) & (n616) & (!n1182)));
	assign n754 = (((!n1009) & (!n527) & (!n638) & (n965)) + ((!n1009) & (!n527) & (n638) & (!n965)) + ((!n1009) & (!n527) & (n638) & (n965)) + ((!n1009) & (n527) & (!n638) & (!n965)) + ((!n1009) & (n527) & (!n638) & (n965)) + ((!n1009) & (n527) & (n638) & (!n965)) + ((!n1009) & (n527) & (n638) & (n965)) + ((n1009) & (!n527) & (!n638) & (!n965)) + ((n1009) & (!n527) & (!n638) & (n965)) + ((n1009) & (!n527) & (n638) & (!n965)) + ((n1009) & (!n527) & (n638) & (n965)) + ((n1009) & (n527) & (!n638) & (!n965)) + ((n1009) & (n527) & (!n638) & (n965)) + ((n1009) & (n527) & (n638) & (!n965)) + ((n1009) & (n527) & (n638) & (n965)));
	assign n755 = (((!n630) & (!n907) & (!i_0_) & (i_8_)) + ((!n630) & (!n907) & (i_0_) & (!i_8_)) + ((!n630) & (!n907) & (i_0_) & (i_8_)) + ((!n630) & (n907) & (!i_0_) & (!i_8_)) + ((!n630) & (n907) & (!i_0_) & (i_8_)) + ((!n630) & (n907) & (i_0_) & (!i_8_)) + ((!n630) & (n907) & (i_0_) & (i_8_)) + ((n630) & (!n907) & (!i_0_) & (!i_8_)) + ((n630) & (!n907) & (!i_0_) & (i_8_)) + ((n630) & (!n907) & (i_0_) & (!i_8_)) + ((n630) & (!n907) & (i_0_) & (i_8_)) + ((n630) & (n907) & (!i_0_) & (!i_8_)) + ((n630) & (n907) & (!i_0_) & (i_8_)) + ((n630) & (n907) & (i_0_) & (!i_8_)) + ((n630) & (n907) & (i_0_) & (i_8_)));
	assign n756 = (((n1198) & (!n641) & (!n241) & (n649)) + ((n1198) & (!n641) & (n241) & (!n649)) + ((n1198) & (!n641) & (n241) & (n649)) + ((n1198) & (n641) & (!n241) & (!n649)) + ((n1198) & (n641) & (!n241) & (n649)) + ((n1198) & (n641) & (n241) & (!n649)) + ((n1198) & (n641) & (n241) & (n649)));
	assign n757 = (((!n608) & (!n1164) & (n1199) & (n1201)) + ((n608) & (!n1164) & (n1199) & (n1201)) + ((n608) & (n1164) & (n1199) & (n1201)));
	assign n758 = (((!i_25_) & (!n448) & (!n740) & (n743)) + ((!i_25_) & (!n448) & (n740) & (n743)) + ((!i_25_) & (n448) & (!n740) & (!n743)) + ((!i_25_) & (n448) & (!n740) & (n743)) + ((!i_25_) & (n448) & (n740) & (!n743)) + ((!i_25_) & (n448) & (n740) & (n743)) + ((i_25_) & (!n448) & (n740) & (n743)) + ((i_25_) & (n448) & (n740) & (!n743)) + ((i_25_) & (n448) & (n740) & (n743)));
	assign n759 = (((!n450) & (n748) & (!n745) & (n1015)) + ((!n450) & (n748) & (n745) & (!n1015)) + ((!n450) & (n748) & (n745) & (n1015)) + ((n450) & (!n748) & (!n745) & (n1015)) + ((n450) & (!n748) & (n745) & (!n1015)) + ((n450) & (!n748) & (n745) & (n1015)) + ((n450) & (n748) & (!n745) & (n1015)) + ((n450) & (n748) & (n745) & (!n1015)) + ((n450) & (n748) & (n745) & (n1015)));
	assign n760 = (((n1202) & (!n884) & (n1172) & (n1203)) + ((n1202) & (n884) & (!n1172) & (!n1203)) + ((n1202) & (n884) & (!n1172) & (n1203)) + ((n1202) & (n884) & (n1172) & (!n1203)) + ((n1202) & (n884) & (n1172) & (n1203)));
	assign n761 = (((!n750) & (!n1033) & (n1204) & (n1205) & (n1206) & (n1207) & (n1208) & (n1210)));
	assign n753 = (((n754) & (n755) & (n756) & (n757) & (n758) & (n759) & (n760) & (n761)));
	assign n763 = (((!i_13_) & (!n735)) + ((!i_13_) & (n735)) + ((i_13_) & (n735)));
	assign n762 = (((!i_12_) & (!i_13_) & (!n453) & (n763)) + ((!i_12_) & (!i_13_) & (n453) & (n763)) + ((!i_12_) & (i_13_) & (n453) & (n763)) + ((i_12_) & (!i_13_) & (!n453) & (!n763)) + ((i_12_) & (!i_13_) & (!n453) & (n763)) + ((i_12_) & (!i_13_) & (n453) & (!n763)) + ((i_12_) & (!i_13_) & (n453) & (n763)) + ((i_12_) & (i_13_) & (n453) & (!n763)) + ((i_12_) & (i_13_) & (n453) & (n763)));
	assign n764 = (((n522) & (n453)));
	assign n765 = (((!i_10_) & (!i_13_) & (!n453) & (n522)) + ((!i_10_) & (!i_13_) & (n453) & (n522)) + ((!i_10_) & (i_13_) & (n453) & (n522)) + ((i_10_) & (!i_13_) & (!n453) & (!n522)) + ((i_10_) & (!i_13_) & (!n453) & (n522)) + ((i_10_) & (!i_13_) & (n453) & (!n522)) + ((i_10_) & (!i_13_) & (n453) & (n522)) + ((i_10_) & (i_13_) & (n453) & (!n522)) + ((i_10_) & (i_13_) & (n453) & (n522)));
	assign n767 = (((!i_3_) & (!i_4_) & (!i_5_)) + ((!i_3_) & (!i_4_) & (i_5_)) + ((!i_3_) & (i_4_) & (!i_5_)) + ((!i_3_) & (i_4_) & (i_5_)) + ((i_3_) & (!i_4_) & (i_5_)) + ((i_3_) & (i_4_) & (!i_5_)) + ((i_3_) & (i_4_) & (i_5_)));
	assign n766 = (((!n586) & (!i_6_) & (n767)) + ((!n586) & (i_6_) & (!n767)) + ((!n586) & (i_6_) & (n767)) + ((n586) & (!i_6_) & (!n767)) + ((n586) & (!i_6_) & (n767)) + ((n586) & (i_6_) & (!n767)) + ((n586) & (i_6_) & (n767)));
	assign n769 = (((!i_4_) & (n373)) + ((i_4_) & (!n373)) + ((i_4_) & (n373)));
	assign n768 = (((!i_2_) & (!i_8_) & (!n769) & (!n951)) + ((!i_2_) & (!i_8_) & (n769) & (!n951)) + ((!i_2_) & (!i_8_) & (n769) & (n951)) + ((!i_2_) & (i_8_) & (!n769) & (!n951)) + ((!i_2_) & (i_8_) & (!n769) & (n951)) + ((!i_2_) & (i_8_) & (n769) & (!n951)) + ((!i_2_) & (i_8_) & (n769) & (n951)));
	assign n771 = (((!i_7_) & (!i_32_) & (i_36_) & (!n769)));
	assign n773 = (((!n765) & (!n768) & (!n771)) + ((!n765) & (!n768) & (n771)) + ((!n765) & (n768) & (n771)));
	assign n777 = (((!i_13_) & (!n575) & (!n766) & (!n769)) + ((!i_13_) & (!n575) & (!n766) & (n769)) + ((!i_13_) & (!n575) & (n766) & (!n769)) + ((!i_13_) & (n575) & (!n766) & (!n769)) + ((!i_13_) & (n575) & (!n766) & (n769)));
	assign n778 = (((!i_32_) & (n951)));
	assign n776 = (((!i_9_) & (!n773) & (n777) & (n778)) + ((!i_9_) & (n773) & (!n777) & (!n778)) + ((!i_9_) & (n773) & (!n777) & (n778)) + ((!i_9_) & (n773) & (n777) & (!n778)) + ((!i_9_) & (n773) & (n777) & (n778)));
	assign n782 = (((!n290) & (!n951) & (n1242) & (!n1241)) + ((!n290) & (!n951) & (n1242) & (n1241)) + ((!n290) & (n951) & (n1242) & (!n1241)) + ((!n290) & (n951) & (n1242) & (n1241)) + ((n290) & (!n951) & (n1242) & (!n1241)) + ((n290) & (!n951) & (n1242) & (n1241)) + ((n290) & (n951) & (n1242) & (n1241)));
	assign n781 = (((!i_31_) & (!n769) & (!n778) & (!n1241)) + ((!i_31_) & (!n769) & (!n778) & (n1241)) + ((!i_31_) & (!n769) & (n778) & (n1241)) + ((!i_31_) & (n769) & (!n778) & (!n1241)) + ((!i_31_) & (n769) & (!n778) & (n1241)) + ((!i_31_) & (n769) & (n778) & (!n1241)) + ((!i_31_) & (n769) & (n778) & (n1241)) + ((i_31_) & (!n769) & (!n778) & (!n1241)) + ((i_31_) & (!n769) & (!n778) & (n1241)) + ((i_31_) & (!n769) & (n778) & (!n1241)) + ((i_31_) & (!n769) & (n778) & (n1241)) + ((i_31_) & (n769) & (!n778) & (!n1241)) + ((i_31_) & (n769) & (!n778) & (n1241)) + ((i_31_) & (n769) & (n778) & (!n1241)) + ((i_31_) & (n769) & (n778) & (n1241)));
	assign n779 = (((!i_29_) & (!n776) & (n782) & (!n781)) + ((!i_29_) & (!n776) & (n782) & (n781)) + ((!i_29_) & (n776) & (n782) & (!n781)) + ((!i_29_) & (n776) & (n782) & (n781)) + ((i_29_) & (!n776) & (n782) & (n781)));
	assign n784 = (((n1261) & (n654)));
	assign n785 = (((n1021) & (n696)));
	assign n783 = (((!i_36_) & (!n784) & (!n785) & (!n951)) + ((!i_36_) & (!n784) & (n785) & (!n951)) + ((!i_36_) & (n784) & (!n785) & (!n951)) + ((!i_36_) & (n784) & (!n785) & (n951)) + ((!i_36_) & (n784) & (n785) & (!n951)) + ((!i_36_) & (n784) & (n785) & (n951)) + ((i_36_) & (!n784) & (n785) & (!n951)) + ((i_36_) & (n784) & (n785) & (!n951)) + ((i_36_) & (n784) & (n785) & (n951)));
	assign n789 = (((!n546) & (n522)) + ((n546) & (!n522)) + ((n546) & (n522)));
	assign n787 = (((!n608) & (!n778) & (n783) & (!n789)) + ((!n608) & (!n778) & (n783) & (n789)) + ((!n608) & (n778) & (n783) & (n789)) + ((n608) & (!n778) & (!n783) & (!n789)) + ((n608) & (!n778) & (!n783) & (n789)) + ((n608) & (!n778) & (n783) & (!n789)) + ((n608) & (!n778) & (n783) & (n789)) + ((n608) & (n778) & (!n783) & (n789)) + ((n608) & (n778) & (n783) & (n789)));
	assign n790 = (((n620) & (n609)));
	assign n792 = (((n607) & (n619)));
	assign n791 = (((!n364) & (!n608) & (n790) & (!n792)) + ((!n364) & (!n608) & (n790) & (n792)) + ((!n364) & (n608) & (!n790) & (!n792)) + ((!n364) & (n608) & (!n790) & (n792)) + ((!n364) & (n608) & (n790) & (!n792)) + ((!n364) & (n608) & (n790) & (n792)) + ((n364) & (!n608) & (n790) & (n792)) + ((n364) & (n608) & (!n790) & (n792)) + ((n364) & (n608) & (n790) & (n792)));
	assign n794 = (((n1259) & (n749)));
	assign n793 = (((!n794) & (n174) & (!n791) & (n243)) + ((!n794) & (n174) & (n791) & (!n243)) + ((!n794) & (n174) & (n791) & (n243)) + ((n794) & (!n174) & (!n791) & (n243)) + ((n794) & (!n174) & (n791) & (!n243)) + ((n794) & (!n174) & (n791) & (n243)) + ((n794) & (n174) & (!n791) & (n243)) + ((n794) & (n174) & (n791) & (!n243)) + ((n794) & (n174) & (n791) & (n243)));
	assign n795 = (((n539) & (!n769)));
	assign n797 = (((!i_9_) & (n769)) + ((i_9_) & (!n769)) + ((i_9_) & (n769)));
	assign n798 = (((n505) & (n763)));
	assign n796 = (((!n229) & (!n531) & (!n797) & (!n798)) + ((!n229) & (!n531) & (!n797) & (n798)) + ((!n229) & (!n531) & (n797) & (!n798)) + ((!n229) & (!n531) & (n797) & (n798)) + ((!n229) & (n531) & (!n797) & (!n798)) + ((!n229) & (n531) & (!n797) & (n798)) + ((!n229) & (n531) & (n797) & (!n798)) + ((!n229) & (n531) & (n797) & (n798)) + ((n229) & (!n531) & (!n797) & (!n798)) + ((n229) & (!n531) & (!n797) & (n798)) + ((n229) & (!n531) & (n797) & (!n798)) + ((n229) & (!n531) & (n797) & (n798)) + ((n229) & (n531) & (!n797) & (n798)) + ((n229) & (n531) & (n797) & (!n798)) + ((n229) & (n531) & (n797) & (n798)));
	assign n801 = (((!i_21_) & (n1003)));
	assign n800 = (((!i_28_) & (n234)));
	assign n799 = (((n13) & (n801) & (!n795) & (n800)) + ((n13) & (n801) & (n795) & (!n800)) + ((n13) & (n801) & (n795) & (n800)));
	assign n802 = (((!i_28_) & (!n785) & (!n796) & (!n1040)) + ((!i_28_) & (!n785) & (n796) & (!n1040)) + ((!i_28_) & (n785) & (!n796) & (!n1040)) + ((i_28_) & (!n785) & (!n796) & (!n1040)) + ((i_28_) & (n785) & (!n796) & (!n1040)));
	assign n806 = (((n367) & (!n1163) & (!n1179)) + ((n367) & (!n1163) & (n1179)) + ((n367) & (n1163) & (!n1179)));
	assign n809 = (((!i_19_) & (!n229) & (!n518) & (!n797)) + ((!i_19_) & (!n229) & (!n518) & (n797)) + ((!i_19_) & (!n229) & (n518) & (!n797)) + ((!i_19_) & (!n229) & (n518) & (n797)) + ((!i_19_) & (n229) & (!n518) & (n797)) + ((!i_19_) & (n229) & (n518) & (!n797)) + ((!i_19_) & (n229) & (n518) & (n797)) + ((i_19_) & (!n229) & (!n518) & (!n797)) + ((i_19_) & (!n229) & (!n518) & (n797)) + ((i_19_) & (!n229) & (n518) & (!n797)) + ((i_19_) & (!n229) & (n518) & (n797)) + ((i_19_) & (n229) & (!n518) & (!n797)) + ((i_19_) & (n229) & (!n518) & (n797)) + ((i_19_) & (n229) & (n518) & (!n797)) + ((i_19_) & (n229) & (n518) & (n797)));
	assign n810 = (((!n767) & (!n640) & (!n98) & (i_18_)) + ((!n767) & (!n640) & (n98) & (!i_18_)) + ((!n767) & (!n640) & (n98) & (i_18_)) + ((!n767) & (n640) & (!n98) & (!i_18_)) + ((!n767) & (n640) & (!n98) & (i_18_)) + ((!n767) & (n640) & (n98) & (!i_18_)) + ((!n767) & (n640) & (n98) & (i_18_)) + ((n767) & (!n640) & (!n98) & (!i_18_)) + ((n767) & (!n640) & (!n98) & (i_18_)) + ((n767) & (!n640) & (n98) & (!i_18_)) + ((n767) & (!n640) & (n98) & (i_18_)) + ((n767) & (n640) & (!n98) & (!i_18_)) + ((n767) & (n640) & (!n98) & (i_18_)) + ((n767) & (n640) & (n98) & (!i_18_)) + ((n767) & (n640) & (n98) & (i_18_)));
	assign n813 = (((!n362) & (!n467)) + ((!n362) & (n467)) + ((n362) & (!n467)));
	assign n812 = (((!i_21_) & (!n833)) + ((i_21_) & (!n833)) + ((i_21_) & (n833)));
	assign n811 = (((n813) & (!n664) & (n812)) + ((n813) & (n664) & (!n812)) + ((n813) & (n664) & (n812)));
	assign n814 = (((!n573) & (!n811) & (!n824)) + ((!n573) & (n811) & (!n824)) + ((n573) & (!n811) & (!n824)));
	assign n818 = (((n467) & (!n644) & (!n659)) + ((n467) & (!n644) & (n659)) + ((n467) & (n644) & (!n659)));
	assign n821 = (((!i_32_) & (n404) & (!n785) & (!n1272)) + ((!i_32_) & (n404) & (!n785) & (n1272)) + ((!i_32_) & (n404) & (n785) & (!n1272)) + ((i_32_) & (n404) & (!n785) & (!n1272)) + ((i_32_) & (n404) & (!n785) & (n1272)));
	assign n826 = (((!n828) & (!n556) & (n444)) + ((!n828) & (n556) & (!n444)) + ((!n828) & (n556) & (n444)) + ((n828) & (!n556) & (!n444)) + ((n828) & (!n556) & (n444)) + ((n828) & (n556) & (!n444)) + ((n828) & (n556) & (n444)));
	assign n824 = (((n1023) & (n695)));
	assign n823 = (((!n653) & (!n821) & (n826) & (n824)) + ((n653) & (!n821) & (n826) & (!n824)) + ((n653) & (!n821) & (n826) & (n824)));
	assign n829 = (((!n215) & (!n367) & (!n1272)) + ((!n215) & (!n367) & (n1272)) + ((!n215) & (n367) & (n1272)) + ((n215) & (!n367) & (!n1272)) + ((n215) & (!n367) & (n1272)) + ((n215) & (n367) & (!n1272)) + ((n215) & (n367) & (n1272)));
	assign n828 = (((n1017) & (n1028)));
	assign n827 = (((!n362) & (!n556) & (n829) & (!n828)) + ((!n362) & (!n556) & (n829) & (n828)) + ((!n362) & (n556) & (n829) & (!n828)) + ((!n362) & (n556) & (n829) & (n828)) + ((n362) & (!n556) & (n829) & (n828)) + ((n362) & (n556) & (n829) & (!n828)) + ((n362) & (n556) & (n829) & (n828)));
	assign n830 = (((!i_7_) & (!n215) & (!n290) & (n785)) + ((!i_7_) & (n215) & (!n290) & (!n785)) + ((!i_7_) & (n215) & (!n290) & (n785)) + ((i_7_) & (!n215) & (!n290) & (n785)) + ((i_7_) & (!n215) & (n290) & (n785)) + ((i_7_) & (n215) & (!n290) & (!n785)) + ((i_7_) & (n215) & (!n290) & (n785)) + ((i_7_) & (n215) & (n290) & (!n785)) + ((i_7_) & (n215) & (n290) & (n785)));
	assign n832 = (((!i_32_) & (i_34_) & (!i_35_)));
	assign n833 = (((!i_23_) & (!i_24_)));
	assign n831 = (((!n243) & (n832) & (n833)));
	assign n834 = (((!n544) & (!n647) & (!n1179)) + ((!n544) & (!n647) & (n1179)) + ((n544) & (!n647) & (!n1179)));
	assign n837 = (((!n570) & (!n642) & (!n659)) + ((!n570) & (!n642) & (n659)) + ((!n570) & (n642) & (!n659)));
	assign n841 = (((!i_29_) & (n253)));
	assign n840 = (((!i_28_) & (!n830) & (!n831) & (n841)) + ((!i_28_) & (!n830) & (n831) & (!n841)) + ((!i_28_) & (!n830) & (n831) & (n841)) + ((!i_28_) & (n830) & (n831) & (!n841)) + ((!i_28_) & (n830) & (n831) & (n841)));
	assign n843 = (((n362) & (!n789) & (!n818) & (n832)) + ((n362) & (!n789) & (n818) & (!n832)) + ((n362) & (!n789) & (n818) & (n832)) + ((n362) & (n789) & (n818) & (!n832)) + ((n362) & (n789) & (n818) & (n832)));
	assign n845 = (((!i_7_) & (!i_32_) & (!n814) & (!n1043)) + ((!i_7_) & (!i_32_) & (n814) & (!n1043)) + ((!i_7_) & (!i_32_) & (n814) & (n1043)) + ((i_7_) & (!i_32_) & (n814) & (!n1043)) + ((i_7_) & (!i_32_) & (n814) & (n1043)));
	assign n847 = (((n10) & (!n799) & (!n802) & (n806)) + ((n10) & (!n799) & (n802) & (!n806)) + ((n10) & (!n799) & (n802) & (n806)) + ((n10) & (n799) & (!n802) & (!n806)) + ((n10) & (n799) & (!n802) & (n806)) + ((n10) & (n799) & (n802) & (!n806)) + ((n10) & (n799) & (n802) & (n806)));
	assign n849 = (((!i_33_) & (!n1004)) + ((!i_33_) & (n1004)) + ((i_33_) & (n1004)));
	assign n848 = (((!n245) & (!n253) & (!n649) & (!n849)) + ((!n245) & (!n253) & (!n649) & (n849)) + ((!n245) & (!n253) & (n649) & (!n849)) + ((!n245) & (!n253) & (n649) & (n849)) + ((!n245) & (n253) & (!n649) & (n849)) + ((!n245) & (n253) & (n649) & (n849)) + ((n245) & (!n253) & (n649) & (!n849)) + ((n245) & (!n253) & (n649) & (n849)) + ((n245) & (n253) & (n649) & (n849)));
	assign n851 = (((n1260) & (n1169)));
	assign n850 = (((n517) & (!i_31_) & (n851)) + ((n517) & (i_31_) & (!n851)) + ((n517) & (i_31_) & (n851)));
	assign n853 = (((n1231) & (!n868) & (!n174) & (n649)) + ((n1231) & (!n868) & (n174) & (!n649)) + ((n1231) & (!n868) & (n174) & (n649)) + ((n1231) & (n868) & (!n174) & (!n649)) + ((n1231) & (n868) & (!n174) & (n649)) + ((n1231) & (n868) & (n174) & (!n649)) + ((n1231) & (n868) & (n174) & (n649)));
	assign n854 = (((!n404) & (!n653) & (!n784) & (n1228)) + ((!n404) & (!n653) & (n784) & (n1228)) + ((!n404) & (n653) & (!n784) & (!n1228)) + ((!n404) & (n653) & (!n784) & (n1228)) + ((!n404) & (n653) & (n784) & (!n1228)) + ((!n404) & (n653) & (n784) & (n1228)) + ((n404) & (!n653) & (n784) & (n1228)) + ((n404) & (n653) & (n784) & (!n1228)) + ((n404) & (n653) & (n784) & (n1228)));
	assign n852 = (((n853) & (n854) & (!n850) & (n444)) + ((n853) & (n854) & (n850) & (!n444)) + ((n853) & (n854) & (n850) & (n444)));
	assign n855 = (((!i_31_) & (n135) & (!n531) & (!n769)) + ((!i_31_) & (n135) & (!n531) & (n769)) + ((!i_31_) & (n135) & (n531) & (n769)) + ((i_31_) & (n135) & (!n531) & (!n769)) + ((i_31_) & (n135) & (!n531) & (n769)) + ((i_31_) & (n135) & (n531) & (!n769)) + ((i_31_) & (n135) & (n531) & (n769)));
	assign n856 = (((!i_8_) & (!n1043)));
	assign n857 = (((n362) & (!n794) & (!n973)));
	assign n859 = (((!i_31_) & (!n811) & (!n856) & (!n1276)) + ((!i_31_) & (!n811) & (n856) & (!n1276)) + ((!i_31_) & (!n811) & (n856) & (n1276)) + ((!i_31_) & (n811) & (n856) & (!n1276)) + ((!i_31_) & (n811) & (n856) & (n1276)));
	assign n861 = (((n10) & (!n350) & (!n517) & (!n1229)) + ((n10) & (!n350) & (n517) & (!n1229)) + ((n10) & (n350) & (!n517) & (!n1229)) + ((n10) & (n350) & (!n517) & (n1229)) + ((n10) & (n350) & (n517) & (!n1229)));
	assign n866 = (((!i_31_) & (!n31) & (!n467) & (!n1004) & (!n1014)) + ((!i_31_) & (!n31) & (!n467) & (!n1004) & (n1014)) + ((!i_31_) & (!n31) & (!n467) & (n1004) & (!n1014)) + ((!i_31_) & (!n31) & (!n467) & (n1004) & (n1014)) + ((!i_31_) & (!n31) & (n467) & (!n1004) & (n1014)) + ((!i_31_) & (!n31) & (n467) & (n1004) & (!n1014)) + ((!i_31_) & (!n31) & (n467) & (n1004) & (n1014)) + ((!i_31_) & (n31) & (!n467) & (!n1004) & (!n1014)) + ((!i_31_) & (n31) & (!n467) & (!n1004) & (n1014)) + ((!i_31_) & (n31) & (!n467) & (n1004) & (!n1014)) + ((!i_31_) & (n31) & (!n467) & (n1004) & (n1014)) + ((!i_31_) & (n31) & (n467) & (!n1004) & (!n1014)) + ((!i_31_) & (n31) & (n467) & (!n1004) & (n1014)) + ((!i_31_) & (n31) & (n467) & (n1004) & (!n1014)) + ((!i_31_) & (n31) & (n467) & (n1004) & (n1014)) + ((i_31_) & (!n31) & (!n467) & (!n1004) & (!n1014)) + ((i_31_) & (!n31) & (!n467) & (!n1004) & (n1014)) + ((i_31_) & (!n31) & (!n467) & (n1004) & (!n1014)) + ((i_31_) & (!n31) & (!n467) & (n1004) & (n1014)) + ((i_31_) & (!n31) & (n467) & (!n1004) & (!n1014)) + ((i_31_) & (!n31) & (n467) & (!n1004) & (n1014)) + ((i_31_) & (!n31) & (n467) & (n1004) & (!n1014)) + ((i_31_) & (!n31) & (n467) & (n1004) & (n1014)) + ((i_31_) & (n31) & (!n467) & (!n1004) & (!n1014)) + ((i_31_) & (n31) & (!n467) & (!n1004) & (n1014)) + ((i_31_) & (n31) & (!n467) & (n1004) & (!n1014)) + ((i_31_) & (n31) & (!n467) & (n1004) & (n1014)) + ((i_31_) & (n31) & (n467) & (!n1004) & (!n1014)) + ((i_31_) & (n31) & (n467) & (!n1004) & (n1014)) + ((i_31_) & (n31) & (n467) & (n1004) & (!n1014)) + ((i_31_) & (n31) & (n467) & (n1004) & (n1014)));
	assign n864 = (((!n681) & (!n797) & (n866) & (!n1044)) + ((!n681) & (!n797) & (n866) & (n1044)) + ((!n681) & (n797) & (n866) & (!n1044)) + ((!n681) & (n797) & (n866) & (n1044)) + ((n681) & (!n797) & (n866) & (!n1044)) + ((n681) & (n797) & (n866) & (!n1044)) + ((n681) & (n797) & (n866) & (n1044)));
	assign n868 = (((n534) & (n704)));
	assign n867 = (((!n10) & (!n170) & (!n868)) + ((!n10) & (!n170) & (n868)) + ((!n10) & (n170) & (!n868)) + ((!n10) & (n170) & (n868)) + ((n10) & (!n170) & (n868)) + ((n10) & (n170) & (!n868)) + ((n10) & (n170) & (n868)));
	assign n870 = (((!i_34_) & (n121) & (!n243)));
	assign n872 = (((!i_14_) & (!i_25_)));
	assign n871 = (((!n497) & (!n872) & (!i_28_) & (i_30_)) + ((!n497) & (!n872) & (i_28_) & (!i_30_)) + ((!n497) & (!n872) & (i_28_) & (i_30_)) + ((!n497) & (n872) & (!i_28_) & (!i_30_)) + ((!n497) & (n872) & (!i_28_) & (i_30_)) + ((!n497) & (n872) & (i_28_) & (!i_30_)) + ((!n497) & (n872) & (i_28_) & (i_30_)) + ((n497) & (!n872) & (!i_28_) & (!i_30_)) + ((n497) & (!n872) & (!i_28_) & (i_30_)) + ((n497) & (!n872) & (i_28_) & (!i_30_)) + ((n497) & (!n872) & (i_28_) & (i_30_)) + ((n497) & (n872) & (!i_28_) & (!i_30_)) + ((n497) & (n872) & (!i_28_) & (i_30_)) + ((n497) & (n872) & (i_28_) & (!i_30_)) + ((n497) & (n872) & (i_28_) & (i_30_)));
	assign n875 = (((!i_24_) & (!n290) & (!n531)) + ((!i_24_) & (!n290) & (n531)) + ((!i_24_) & (n290) & (!n531)) + ((i_24_) & (!n290) & (!n531)) + ((i_24_) & (!n290) & (n531)) + ((i_24_) & (n290) & (!n531)) + ((i_24_) & (n290) & (n531)));
	assign n874 = (((n479) & (!n688)));
	assign n873 = (((!i_29_) & (!n649) & (n875) & (!n874)) + ((!i_29_) & (!n649) & (n875) & (n874)) + ((!i_29_) & (n649) & (n875) & (!n874)) + ((!i_29_) & (n649) & (n875) & (n874)) + ((i_29_) & (!n649) & (n875) & (n874)) + ((i_29_) & (n649) & (n875) & (!n874)) + ((i_29_) & (n649) & (n875) & (n874)));
	assign n880 = (((n833) & (i_21_)));
	assign n876 = (((!n723) & (!n871) & (n880) & (!n1038)) + ((!n723) & (!n871) & (n880) & (n1038)) + ((!n723) & (n871) & (n880) & (!n1038)) + ((n723) & (!n871) & (n880) & (!n1038)) + ((n723) & (!n871) & (n880) & (n1038)));
	assign n882 = (((!n10) & (!n238) & (n649) & (!n995)) + ((!n10) & (!n238) & (n649) & (n995)) + ((!n10) & (n238) & (!n649) & (!n995)) + ((!n10) & (n238) & (!n649) & (n995)) + ((!n10) & (n238) & (n649) & (!n995)) + ((!n10) & (n238) & (n649) & (n995)) + ((n10) & (!n238) & (n649) & (n995)) + ((n10) & (n238) & (!n649) & (n995)) + ((n10) & (n238) & (n649) & (n995)));
	assign n881 = (((!n211) & (!n362) & (n882)) + ((n211) & (!n362) & (n882)) + ((n211) & (n362) & (n882)));
	assign n884 = (((!i_23_) & (n1004)) + ((i_23_) & (!n1004)) + ((i_23_) & (n1004)));
	assign n883 = (((!n884) & (n211) & (!n572) & (n236)) + ((!n884) & (n211) & (n572) & (!n236)) + ((!n884) & (n211) & (n572) & (n236)) + ((n884) & (!n211) & (!n572) & (n236)) + ((n884) & (!n211) & (n572) & (!n236)) + ((n884) & (!n211) & (n572) & (n236)) + ((n884) & (n211) & (!n572) & (n236)) + ((n884) & (n211) & (n572) & (!n236)) + ((n884) & (n211) & (n572) & (n236)));
	assign n886 = (((!i_21_) & (!n883) & (!n1006)) + ((!i_21_) & (!n883) & (n1006)) + ((!i_21_) & (n883) & (!n1006)) + ((!i_21_) & (n883) & (n1006)) + ((i_21_) & (!n883) & (n1006)) + ((i_21_) & (n883) & (!n1006)) + ((i_21_) & (n883) & (n1006)));
	assign n885 = (((n886) & (!n881) & (n556)) + ((n886) & (n881) & (!n556)) + ((n886) & (n881) & (n556)));
	assign n888 = (((!i_11_) & (n1036)) + ((i_11_) & (!n1036)) + ((i_11_) & (n1036)));
	assign n889 = (((!i_3_) & (!n1036)) + ((!i_3_) & (n1036)) + ((i_3_) & (n1036)));
	assign n887 = (((!i_19_) & (n888) & (!i_18_) & (n889)) + ((!i_19_) & (n888) & (i_18_) & (!n889)) + ((!i_19_) & (n888) & (i_18_) & (n889)) + ((i_19_) & (!n888) & (!i_18_) & (n889)) + ((i_19_) & (!n888) & (i_18_) & (!n889)) + ((i_19_) & (!n888) & (i_18_) & (n889)) + ((i_19_) & (n888) & (!i_18_) & (n889)) + ((i_19_) & (n888) & (i_18_) & (!n889)) + ((i_19_) & (n888) & (i_18_) & (n889)));
	assign n891 = (((i_21_) & (!i_23_)));
	assign n890 = (((i_25_) & (!n849) & (n891)));
	assign n892 = (((n290) & (n531) & (i_22_)));
	assign n893 = (((!n479) & (!n672) & (!n673) & (n890)) + ((!n479) & (!n672) & (n673) & (n890)) + ((!n479) & (n672) & (!n673) & (n890)) + ((!n479) & (n672) & (n673) & (!n890)) + ((!n479) & (n672) & (n673) & (n890)));
	assign n895 = (((!i_18_) & (!n81) & (n767)) + ((!i_18_) & (n81) & (!n767)) + ((!i_18_) & (n81) & (n767)) + ((i_18_) & (!n81) & (!n767)) + ((i_18_) & (!n81) & (n767)) + ((i_18_) & (n81) & (!n767)) + ((i_18_) & (n81) & (n767)));
	assign n894 = (((!i_7_) & (!n19) & (!n797) & (n895)) + ((!i_7_) & (!n19) & (n797) & (n895)) + ((!i_7_) & (n19) & (n797) & (n895)) + ((i_7_) & (!n19) & (!n797) & (n895)) + ((i_7_) & (!n19) & (n797) & (n895)) + ((i_7_) & (n19) & (!n797) & (n895)) + ((i_7_) & (n19) & (n797) & (n895)));
	assign n897 = (((!i_2_) & (!i_3_) & (!i_9_)) + ((!i_2_) & (!i_3_) & (i_9_)) + ((!i_2_) & (i_3_) & (!i_9_)) + ((!i_2_) & (i_3_) & (i_9_)) + ((i_2_) & (!i_3_) & (!i_9_)) + ((i_2_) & (!i_3_) & (i_9_)) + ((i_2_) & (i_3_) & (i_9_)));
	assign n896 = (((!n84) & (!n767) & (n897) & (!n951)) + ((!n84) & (n767) & (n897) & (!n951)) + ((!n84) & (n767) & (n897) & (n951)) + ((n84) & (!n767) & (n897) & (!n951)) + ((n84) & (!n767) & (n897) & (n951)) + ((n84) & (n767) & (n897) & (!n951)) + ((n84) & (n767) & (n897) & (n951)));
	assign n898 = (((!i_9_) & (n19) & (!n768)));
	assign n899 = (((!i_18_) & (n531) & (!n896) & (!n898)) + ((!i_18_) & (n531) & (!n896) & (n898)) + ((!i_18_) & (n531) & (n896) & (n898)) + ((i_18_) & (n531) & (!n896) & (n898)) + ((i_18_) & (n531) & (n896) & (n898)));
	assign n901 = (((!i_36_) & (!n539) & (!n894) & (!n899)) + ((!i_36_) & (!n539) & (n894) & (!n899)) + ((!i_36_) & (n539) & (!n894) & (!n899)) + ((!i_36_) & (n539) & (n894) & (!n899)) + ((i_36_) & (!n539) & (!n894) & (!n899)) + ((i_36_) & (!n539) & (n894) & (!n899)) + ((i_36_) & (n539) & (n894) & (!n899)));
	assign n904 = (((!i_31_) & (!n334) & (!n692) & (!n1279)) + ((!i_31_) & (n334) & (!n692) & (!n1279)) + ((!i_31_) & (n334) & (n692) & (!n1279)) + ((i_31_) & (!n334) & (!n692) & (!n1279)) + ((i_31_) & (!n334) & (n692) & (!n1279)) + ((i_31_) & (n334) & (!n692) & (!n1279)) + ((i_31_) & (n334) & (n692) & (!n1279)));
	assign n907 = (((!n467) & (!n1005)) + ((!n467) & (n1005)) + ((n467) & (n1005)));
	assign n906 = (((!n681) & (!n769) & (n907)) + ((!n681) & (n769) & (n907)) + ((n681) & (n769) & (n907)));
	assign n909 = (((!n192) & (!n608) & (n664)) + ((!n192) & (n608) & (!n664)) + ((!n192) & (n608) & (n664)) + ((n192) & (!n608) & (!n664)) + ((n192) & (!n608) & (n664)) + ((n192) & (n608) & (!n664)) + ((n192) & (n608) & (n664)));
	assign n908 = (((!n11) & (!n215) & (!n334) & (n909)) + ((!n11) & (!n215) & (n334) & (n909)) + ((!n11) & (n215) & (!n334) & (n909)) + ((!n11) & (n215) & (n334) & (n909)) + ((n11) & (!n215) & (n334) & (n909)) + ((n11) & (n215) & (!n334) & (n909)) + ((n11) & (n215) & (n334) & (n909)));
	assign n911 = (((!i_34_) & (!i_36_) & (!n234)) + ((!i_34_) & (!i_36_) & (n234)) + ((!i_34_) & (i_36_) & (!n234)) + ((!i_34_) & (i_36_) & (n234)) + ((i_34_) & (!i_36_) & (!n234)) + ((i_34_) & (!i_36_) & (n234)) + ((i_34_) & (i_36_) & (!n234)));
	assign n910 = (((!i_36_) & (!n404) & (!n908) & (!n911)) + ((!i_36_) & (!n404) & (!n908) & (n911)) + ((!i_36_) & (!n404) & (n908) & (!n911)) + ((!i_36_) & (!n404) & (n908) & (n911)) + ((!i_36_) & (n404) & (!n908) & (n911)) + ((!i_36_) & (n404) & (n908) & (n911)) + ((i_36_) & (!n404) & (n908) & (!n911)) + ((i_36_) & (!n404) & (n908) & (n911)) + ((i_36_) & (n404) & (n908) & (n911)));
	assign n912 = (((!i_2_) & (!n135) & (!n778)) + ((!i_2_) & (n135) & (!n778)) + ((!i_2_) & (n135) & (n778)) + ((i_2_) & (!n135) & (!n778)) + ((i_2_) & (!n135) & (n778)) + ((i_2_) & (n135) & (!n778)) + ((i_2_) & (n135) & (n778)));
	assign n916 = (((!n9) & (!n229) & (!n556) & (!n1281)) + ((!n9) & (!n229) & (n556) & (!n1281)) + ((!n9) & (n229) & (!n556) & (!n1281)) + ((!n9) & (n229) & (n556) & (!n1281)) + ((n9) & (!n229) & (!n556) & (!n1281)) + ((n9) & (!n229) & (n556) & (!n1281)) + ((n9) & (n229) & (n556) & (!n1281)));
	assign n914 = (((!i_7_) & (n910) & (!n1040) & (!n1216)) + ((!i_7_) & (n910) & (n1040) & (!n1216)) + ((!i_7_) & (n910) & (n1040) & (n1216)) + ((i_7_) & (!n910) & (!n1040) & (!n1216)) + ((i_7_) & (!n910) & (n1040) & (!n1216)) + ((i_7_) & (!n910) & (n1040) & (n1216)) + ((i_7_) & (n910) & (!n1040) & (!n1216)) + ((i_7_) & (n910) & (n1040) & (!n1216)) + ((i_7_) & (n910) & (n1040) & (n1216)));
	assign n915 = (((!i_21_) & (!n883) & (!n931) & (n1257)) + ((!i_21_) & (!n883) & (n931) & (n1257)) + ((!i_21_) & (n883) & (!n931) & (n1257)) + ((!i_21_) & (n883) & (n931) & (n1257)) + ((i_21_) & (!n883) & (n931) & (n1257)) + ((i_21_) & (n883) & (!n931) & (n1257)) + ((i_21_) & (n883) & (n931) & (n1257)));
	assign n913 = (((n916) & (!i_16_) & (n914) & (n915)) + ((n916) & (i_16_) & (!n914) & (!n915)) + ((n916) & (i_16_) & (!n914) & (n915)) + ((n916) & (i_16_) & (n914) & (!n915)) + ((n916) & (i_16_) & (n914) & (n915)));
	assign n917 = (((!n548) & (n888) & (!n547) & (n889)) + ((!n548) & (n888) & (n547) & (!n889)) + ((!n548) & (n888) & (n547) & (n889)) + ((n548) & (!n888) & (!n547) & (n889)) + ((n548) & (!n888) & (n547) & (!n889)) + ((n548) & (!n888) & (n547) & (n889)) + ((n548) & (n888) & (!n547) & (n889)) + ((n548) & (n888) & (n547) & (!n889)) + ((n548) & (n888) & (n547) & (n889)));
	assign n919 = (((!n722) & (!n887) & (!n891)) + ((!n722) & (n887) & (!n891)) + ((!n722) & (n887) & (n891)) + ((n722) & (!n887) & (!n891)) + ((n722) & (!n887) & (n891)) + ((n722) & (n887) & (!n891)) + ((n722) & (n887) & (n891)));
	assign n918 = (((n919) & (!n725) & (n917)) + ((n919) & (n725) & (!n917)) + ((n919) & (n725) & (n917)));
	assign n920 = (((!i_16_) & (!i_17_) & (n216) & (!n363)) + ((!i_16_) & (i_17_) & (!n216) & (!n363)) + ((!i_16_) & (i_17_) & (n216) & (!n363)) + ((i_16_) & (!i_17_) & (n216) & (!n363)) + ((i_16_) & (!i_17_) & (n216) & (n363)) + ((i_16_) & (i_17_) & (!n216) & (!n363)) + ((i_16_) & (i_17_) & (!n216) & (n363)) + ((i_16_) & (i_17_) & (n216) & (!n363)) + ((i_16_) & (i_17_) & (n216) & (n363)));
	assign n922 = (((!n497) & (n741)) + ((n497) & (!n741)) + ((n497) & (n741)));
	assign n921 = (((!i_21_) & (!n407) & (!n737) & (n922)) + ((!i_21_) & (!n407) & (n737) & (n922)) + ((i_21_) & (!n407) & (n737) & (n922)));
	assign n926 = (((!n791) & (!n1039) & (!i_31_) & (i_30_)) + ((!n791) & (!n1039) & (i_31_) & (!i_30_)) + ((!n791) & (!n1039) & (i_31_) & (i_30_)) + ((!n791) & (n1039) & (!i_31_) & (!i_30_)) + ((!n791) & (n1039) & (!i_31_) & (i_30_)) + ((!n791) & (n1039) & (i_31_) & (!i_30_)) + ((!n791) & (n1039) & (i_31_) & (i_30_)) + ((n791) & (!n1039) & (!i_31_) & (!i_30_)) + ((n791) & (!n1039) & (!i_31_) & (i_30_)) + ((n791) & (!n1039) & (i_31_) & (!i_30_)) + ((n791) & (!n1039) & (i_31_) & (i_30_)) + ((n791) & (n1039) & (!i_31_) & (!i_30_)) + ((n791) & (n1039) & (!i_31_) & (i_30_)) + ((n791) & (n1039) & (i_31_) & (!i_30_)) + ((n791) & (n1039) & (i_31_) & (i_30_)));
	assign n924 = (((!n13) & (!n364) & (!n911) & (n926)) + ((!n13) & (!n364) & (n911) & (n926)) + ((!n13) & (n364) & (!n911) & (n926)) + ((!n13) & (n364) & (n911) & (n926)) + ((n13) & (!n364) & (!n911) & (n926)) + ((n13) & (!n364) & (n911) & (n926)) + ((n13) & (n364) & (n911) & (n926)));
	assign n927 = (((!i_31_) & (!n467) & (!n573) & (!n723)) + ((!i_31_) & (!n467) & (!n573) & (n723)) + ((!i_31_) & (!n467) & (n573) & (!n723)) + ((!i_31_) & (!n467) & (n573) & (n723)) + ((!i_31_) & (n467) & (!n573) & (n723)) + ((!i_31_) & (n467) & (n573) & (n723)) + ((i_31_) & (!n467) & (n573) & (!n723)) + ((i_31_) & (!n467) & (n573) & (n723)) + ((i_31_) & (n467) & (n573) & (n723)));
	assign n931 = (((!i_12_) & (n1035)) + ((i_12_) & (!n1035)) + ((i_12_) & (n1035)));
	assign n929 = (((!n9) & (!n559) & (!n881) & (n931)) + ((!n9) & (!n559) & (n881) & (!n931)) + ((!n9) & (!n559) & (n881) & (n931)) + ((!n9) & (n559) & (!n881) & (n931)) + ((!n9) & (n559) & (n881) & (!n931)) + ((!n9) & (n559) & (n881) & (n931)) + ((n9) & (n559) & (!n881) & (n931)) + ((n9) & (n559) & (n881) & (!n931)) + ((n9) & (n559) & (n881) & (n931)));
	assign n939 = (((!i_20_) & (!i_21_) & (!n904) & (!n1280)) + ((!i_20_) & (!i_21_) & (n904) & (!n1280)) + ((i_20_) & (!i_21_) & (!n904) & (!n1280)) + ((i_20_) & (!i_21_) & (!n904) & (n1280)) + ((i_20_) & (!i_21_) & (n904) & (!n1280)));
	assign n942 = (((n253) & (!n892) & (!n893) & (!n1223)) + ((n253) & (!n892) & (n893) & (!n1223)) + ((n253) & (!n892) & (n893) & (n1223)) + ((n253) & (n892) & (!n893) & (!n1223)) + ((n253) & (n892) & (!n893) & (n1223)) + ((n253) & (n892) & (n893) & (!n1223)) + ((n253) & (n892) & (n893) & (n1223)));
	assign n944 = (((i_34_) & (!n496) & (!n876) & (!n1224)) + ((i_34_) & (!n496) & (!n876) & (n1224)) + ((i_34_) & (!n496) & (n876) & (!n1224)) + ((i_34_) & (!n496) & (n876) & (n1224)) + ((i_34_) & (n496) & (!n876) & (!n1224)) + ((i_34_) & (n496) & (n876) & (!n1224)) + ((i_34_) & (n496) & (n876) & (n1224)));
	assign n947 = (((n778) & (!n867) & (!n870) & (!n1227)) + ((n778) & (!n867) & (!n870) & (n1227)) + ((n778) & (!n867) & (n870) & (!n1227)) + ((n778) & (!n867) & (n870) & (n1227)) + ((n778) & (n867) & (!n870) & (!n1227)) + ((n778) & (n867) & (n870) & (!n1227)) + ((n778) & (n867) & (n870) & (n1227)));
	assign n951 = (((!i_35_) & (i_36_)));
	assign n950 = (((n951) & (!n857) & (!n859) & (n861)) + ((n951) & (!n857) & (n859) & (!n861)) + ((n951) & (!n857) & (n859) & (n861)) + ((n951) & (n857) & (!n859) & (!n861)) + ((n951) & (n857) & (!n859) & (n861)) + ((n951) & (n857) & (n859) & (!n861)) + ((n951) & (n857) & (n859) & (n861)));
	assign n953 = (((!i_12_) & (n735)) + ((i_12_) & (!n735)) + ((i_12_) & (n735)));
	assign n954 = (((!i_21_) & (i_22_)) + ((i_21_) & (!i_22_)) + ((i_21_) & (i_22_)));
	assign n957 = (((!i_16_) & (!i_27_)));
	assign n960 = (((!i_23_) & (i_17_)) + ((i_23_) & (!i_17_)) + ((i_23_) & (i_17_)));
	assign n961 = (((!i_2_) & (i_4_)) + ((i_2_) & (!i_4_)) + ((i_2_) & (i_4_)));
	assign n962 = (((!i_9_) & (!n373)) + ((!i_9_) & (n373)) + ((i_9_) & (n373)));
	assign n963 = (((!i_28_) & (i_26_)) + ((i_28_) & (!i_26_)) + ((i_28_) & (i_26_)));
	assign n964 = (((!i_8_) & (!i_9_)) + ((i_8_) & (!i_9_)) + ((i_8_) & (i_9_)));
	assign n965 = (((!i_8_) & (n373)) + ((i_8_) & (!n373)) + ((i_8_) & (n373)));
	assign n966 = (((!i_2_) & (i_3_)) + ((i_2_) & (!i_3_)) + ((i_2_) & (i_3_)));
	assign n968 = (((!i_33_) & (!n234)) + ((i_33_) & (!n234)) + ((i_33_) & (n234)));
	assign n969 = (((!i_9_) & (!n966)) + ((!i_9_) & (n966)) + ((i_9_) & (n966)));
	assign n970 = (((!i_33_) & (i_32_)) + ((i_33_) & (!i_32_)) + ((i_33_) & (i_32_)));
	assign n972 = (((!i_31_) & (n970)) + ((i_31_) & (!n970)) + ((i_31_) & (n970)));
	assign n973 = (((!i_34_) & (!n685)) + ((!i_34_) & (n685)) + ((i_34_) & (n685)));
	assign n974 = (((!i_30_) & (i_29_)) + ((i_30_) & (!i_29_)) + ((i_30_) & (i_29_)));
	assign n975 = (((!i_8_) & (n372)) + ((i_8_) & (!n372)) + ((i_8_) & (n372)));
	assign n977 = (((!i_4_) & (n966)) + ((i_4_) & (!n966)) + ((i_4_) & (n966)));
	assign n978 = (((!i_29_) & (!i_34_)) + ((i_29_) & (!i_34_)) + ((i_29_) & (i_34_)));
	assign n979 = (((!i_9_) & (!n23)) + ((!i_9_) & (n23)) + ((i_9_) & (!n23)));
	assign n983 = (((!i_3_) & (!n961)) + ((!i_3_) & (n961)) + ((i_3_) & (n961)));
	assign n984 = (((!n983) & (n595)) + ((n983) & (!n595)) + ((n983) & (n595)));
	assign n985 = (((!i_9_) & (n984)) + ((i_9_) & (!n984)) + ((i_9_) & (n984)));
	assign n986 = (((!n371) & (n98)) + ((n371) & (!n98)) + ((n371) & (n98)));
	assign n987 = (((!i_3_) & (!i_7_) & (!i_10_)) + ((!i_3_) & (i_7_) & (!i_10_)) + ((!i_3_) & (i_7_) & (i_10_)) + ((i_3_) & (!i_7_) & (!i_10_)) + ((i_3_) & (!i_7_) & (i_10_)) + ((i_3_) & (i_7_) & (!i_10_)) + ((i_3_) & (i_7_) & (i_10_)));
	assign n988 = (((!i_33_) & (!i_34_) & (!i_35_)) + ((!i_33_) & (!i_34_) & (i_35_)) + ((!i_33_) & (i_34_) & (i_35_)) + ((i_33_) & (!i_34_) & (!i_35_)) + ((i_33_) & (!i_34_) & (i_35_)) + ((i_33_) & (i_34_) & (!i_35_)) + ((i_33_) & (i_34_) & (i_35_)));
	assign n989 = (((!i_9_) & (i_6_)) + ((i_9_) & (!i_6_)) + ((i_9_) & (i_6_)));
	assign n990 = (((!n965) & (n983)) + ((n965) & (!n983)) + ((n965) & (n983)));
	assign n991 = (((!i_11_) & (n989)) + ((i_11_) & (!n989)) + ((i_11_) & (n989)));
	assign n992 = (((!i_7_) & (n372)) + ((i_7_) & (!n372)) + ((i_7_) & (n372)));
	assign n993 = (((!n11) & (!n833)) + ((!n11) & (n833)) + ((n11) & (!n833)));
	assign n994 = (((!n394) & (!n974)) + ((!n394) & (n974)) + ((n394) & (n974)));
	assign n995 = (((!i_28_) & (!i_31_)) + ((i_28_) & (!i_31_)) + ((i_28_) & (i_31_)));
	assign n996 = (((!i_7_) & (!i_28_) & (n192)) + ((!i_7_) & (i_28_) & (!n192)) + ((!i_7_) & (i_28_) & (n192)) + ((i_7_) & (!i_28_) & (!n192)) + ((i_7_) & (!i_28_) & (n192)) + ((i_7_) & (i_28_) & (!n192)) + ((i_7_) & (i_28_) & (n192)));
	assign n997 = (((!i_8_) & (n966)) + ((i_8_) & (!n966)) + ((i_8_) & (n966)));
	assign n998 = (((!i_22_) & (!n531) & (!n874) & (!n891)) + ((!i_22_) & (!n531) & (!n874) & (n891)) + ((!i_22_) & (!n531) & (n874) & (!n891)) + ((!i_22_) & (!n531) & (n874) & (n891)) + ((!i_22_) & (n531) & (!n874) & (!n891)) + ((!i_22_) & (n531) & (n874) & (!n891)) + ((!i_22_) & (n531) & (n874) & (n891)) + ((i_22_) & (!n531) & (!n874) & (!n891)) + ((i_22_) & (!n531) & (!n874) & (n891)) + ((i_22_) & (!n531) & (n874) & (!n891)) + ((i_22_) & (!n531) & (n874) & (n891)) + ((i_22_) & (n531) & (!n874) & (!n891)) + ((i_22_) & (n531) & (!n874) & (n891)) + ((i_22_) & (n531) & (n874) & (!n891)) + ((i_22_) & (n531) & (n874) & (n891)));
	assign n1000 = (((!i_12_) & (!n962) & (n977)) + ((!i_12_) & (n962) & (!n977)) + ((!i_12_) & (n962) & (n977)) + ((i_12_) & (!n962) & (!n977)) + ((i_12_) & (!n962) & (n977)) + ((i_12_) & (n962) & (!n977)) + ((i_12_) & (n962) & (n977)));
	assign n1001 = (((!i_2_) & (!i_7_) & (!i_38_)) + ((!i_2_) & (i_7_) & (!i_38_)) + ((!i_2_) & (i_7_) & (i_38_)) + ((i_2_) & (!i_7_) & (!i_38_)) + ((i_2_) & (!i_7_) & (i_38_)) + ((i_2_) & (i_7_) & (!i_38_)) + ((i_2_) & (i_7_) & (i_38_)));
	assign n1002 = (((!n30) & (n31)) + ((n30) & (!n31)) + ((n30) & (n31)));
	assign n1003 = (((!i_16_) & (!i_23_)));
	assign n1004 = (((!i_27_) & (i_28_)) + ((i_27_) & (!i_28_)) + ((i_27_) & (i_28_)));
	assign n1005 = (((!i_30_) & (n1004)) + ((i_30_) & (!n1004)) + ((i_30_) & (n1004)));
	assign n1006 = (((!i_16_) & (i_17_)) + ((i_16_) & (!i_17_)) + ((i_16_) & (i_17_)));
	assign n1007 = (((!i_0_) & (i_4_)) + ((i_0_) & (!i_4_)) + ((i_0_) & (i_4_)));
	assign n1008 = (((!i_17_) & (!i_20_) & (!n681)) + ((!i_17_) & (i_20_) & (!n681)) + ((!i_17_) & (i_20_) & (n681)) + ((i_17_) & (!i_20_) & (!n681)) + ((i_17_) & (!i_20_) & (n681)) + ((i_17_) & (i_20_) & (!n681)) + ((i_17_) & (i_20_) & (n681)));
	assign n1009 = (((!i_18_) & (n1008)) + ((i_18_) & (!n1008)) + ((i_18_) & (n1008)));
	assign n1010 = (((!i_19_) & (n1006)) + ((i_19_) & (!n1006)) + ((i_19_) & (n1006)));
	assign n1011 = (((!i_12_) & (n734)) + ((i_12_) & (!n734)) + ((i_12_) & (n734)));
	assign n1012 = (((!n371) & (n992)) + ((n371) & (!n992)) + ((n371) & (n992)));
	assign n1013 = (((!i_18_) & (n960)) + ((i_18_) & (!n960)) + ((i_18_) & (n960)));
	assign n1014 = (((!n373) & (n374)) + ((n373) & (!n374)) + ((n373) & (n374)));
	assign n1015 = (((!i_5_) & (n1007)) + ((i_5_) & (!n1007)) + ((i_5_) & (n1007)));
	assign n1016 = (((!n98) & (n1015)) + ((n98) & (!n1015)) + ((n98) & (n1015)));
	assign n1017 = (((!i_13_) & (!i_14_) & (!n70)) + ((!i_13_) & (!i_14_) & (n70)) + ((!i_13_) & (i_14_) & (!n70)) + ((!i_13_) & (i_14_) & (n70)) + ((i_13_) & (!i_14_) & (n70)) + ((i_13_) & (i_14_) & (!n70)) + ((i_13_) & (i_14_) & (n70)));
	assign n1018 = (((!n371) & (n975)) + ((n371) & (!n975)) + ((n371) & (n975)));
	assign n1019 = (((!i_23_) & (n735)) + ((i_23_) & (!n735)) + ((i_23_) & (n735)));
	assign n1020 = (((!i_13_) & (!n989)) + ((!i_13_) & (n989)) + ((i_13_) & (n989)));
	assign n1021 = (((!n96) & (n620)) + ((n96) & (!n620)) + ((n96) & (n620)));
	assign n1022 = (((!n63) & (n453)) + ((n63) & (!n453)) + ((n63) & (n453)));
	assign n1023 = (((!n96) & (n453)) + ((n96) & (!n453)) + ((n96) & (n453)));
	assign n1024 = (((!i_23_) & (!i_27_)));
	assign n1025 = (((!i_25_) & (!n1004)) + ((!i_25_) & (n1004)) + ((i_25_) & (n1004)));
	assign n1026 = (((!i_20_) & (!n833)) + ((!i_20_) & (n833)) + ((i_20_) & (!n833)));
	assign n1027 = (((!i_20_) & (!n833)) + ((i_20_) & (!n833)) + ((i_20_) & (n833)));
	assign n1028 = (((!i_13_) & (!i_10_) & (n70)) + ((!i_13_) & (i_10_) & (!n70)) + ((!i_13_) & (i_10_) & (n70)) + ((i_13_) & (!i_10_) & (!n70)) + ((i_13_) & (!i_10_) & (n70)) + ((i_13_) & (i_10_) & (!n70)) + ((i_13_) & (i_10_) & (n70)));
	assign n1029 = (((!n66) & (n505)) + ((n66) & (!n505)) + ((n66) & (n505)));
	assign n1030 = (((!i_14_) & (i_12_)) + ((i_14_) & (!i_12_)) + ((i_14_) & (i_12_)));
	assign n1033 = (((!n679) & (!n683) & (!n686) & (!n691)) + ((!n679) & (!n683) & (!n686) & (n691)) + ((!n679) & (!n683) & (n686) & (!n691)) + ((!n679) & (!n683) & (n686) & (n691)) + ((!n679) & (n683) & (!n686) & (n691)) + ((!n679) & (n683) & (n686) & (!n691)) + ((!n679) & (n683) & (n686) & (n691)) + ((n679) & (!n683) & (!n686) & (!n691)) + ((n679) & (!n683) & (!n686) & (n691)) + ((n679) & (!n683) & (n686) & (!n691)) + ((n679) & (!n683) & (n686) & (n691)) + ((n679) & (n683) & (!n686) & (!n691)) + ((n679) & (n683) & (!n686) & (n691)) + ((n679) & (n683) & (n686) & (!n691)) + ((n679) & (n683) & (n686) & (n691)));
	assign n1035 = (((!i_7_) & (!i_9_)) + ((!i_7_) & (i_9_)) + ((i_7_) & (i_9_)));
	assign n1036 = (((!i_7_) & (!i_10_)) + ((!i_7_) & (i_10_)) + ((i_7_) & (!i_10_)));
	assign n1038 = (((!n762) & (n1036)) + ((n762) & (!n1036)) + ((n762) & (n1036)));
	assign n1039 = (((!i_34_) & (!n951)) + ((!i_34_) & (n951)) + ((i_34_) & (!n951)));
	assign n1040 = (((!i_21_) & (n960)) + ((i_21_) & (!n960)) + ((i_21_) & (n960)));
	assign n1041 = (((!i_20_) & (!i_21_) & (!i_23_)) + ((!i_20_) & (!i_21_) & (i_23_)) + ((!i_20_) & (i_21_) & (!i_23_)) + ((!i_20_) & (i_21_) & (i_23_)) + ((i_20_) & (!i_21_) & (i_23_)) + ((i_20_) & (i_21_) & (!i_23_)) + ((i_20_) & (i_21_) & (i_23_)));
	assign n1042 = (((!i_21_) & (n1006)) + ((i_21_) & (!n1006)) + ((i_21_) & (n1006)));
	assign n1043 = (((!n907) & (!n1042) & (!i_2_) & (n31)) + ((!n907) & (!n1042) & (i_2_) & (!n31)) + ((!n907) & (!n1042) & (i_2_) & (n31)) + ((!n907) & (n1042) & (!i_2_) & (!n31)) + ((!n907) & (n1042) & (!i_2_) & (n31)) + ((!n907) & (n1042) & (i_2_) & (!n31)) + ((!n907) & (n1042) & (i_2_) & (n31)) + ((n907) & (!n1042) & (!i_2_) & (!n31)) + ((n907) & (!n1042) & (!i_2_) & (n31)) + ((n907) & (!n1042) & (i_2_) & (!n31)) + ((n907) & (!n1042) & (i_2_) & (n31)) + ((n907) & (n1042) & (!i_2_) & (!n31)) + ((n907) & (n1042) & (!i_2_) & (n31)) + ((n907) & (n1042) & (i_2_) & (!n31)) + ((n907) & (n1042) & (i_2_) & (n31)));
	assign n1044 = (((!i_10_) & (!i_13_) & (!i_14_)) + ((!i_10_) & (!i_13_) & (i_14_)) + ((!i_10_) & (i_13_) & (!i_14_)) + ((i_10_) & (i_13_) & (!i_14_)));
	assign n1045 = (((!n170) & (n376) & (!n86) & (n174)) + ((!n170) & (n376) & (n86) & (!n174)) + ((!n170) & (n376) & (n86) & (n174)) + ((n170) & (!n376) & (!n86) & (n174)) + ((n170) & (!n376) & (n86) & (!n174)) + ((n170) & (!n376) & (n86) & (n174)) + ((n170) & (n376) & (!n86) & (n174)) + ((n170) & (n376) & (n86) & (!n174)) + ((n170) & (n376) & (n86) & (n174)));
	assign n1046 = (((!n195) & (!n313) & (n972) & (!n973)) + ((!n195) & (!n313) & (n972) & (n973)) + ((!n195) & (n313) & (n972) & (n973)) + ((n195) & (!n313) & (!n972) & (!n973)) + ((n195) & (!n313) & (!n972) & (n973)) + ((n195) & (!n313) & (n972) & (!n973)) + ((n195) & (!n313) & (n972) & (n973)) + ((n195) & (n313) & (!n972) & (n973)) + ((n195) & (n313) & (n972) & (n973)));
	assign n1047 = (((!n15) & (!n38) & (!n72) & (n261)) + ((!n15) & (!n38) & (n72) & (n261)) + ((!n15) & (n38) & (!n72) & (!n261)) + ((!n15) & (n38) & (!n72) & (n261)) + ((!n15) & (n38) & (n72) & (!n261)) + ((!n15) & (n38) & (n72) & (n261)) + ((n15) & (!n38) & (n72) & (n261)) + ((n15) & (n38) & (n72) & (!n261)) + ((n15) & (n38) & (n72) & (n261)));
	assign n1048 = (((!n23) & (!n64) & (!n63) & (n979)) + ((!n23) & (!n64) & (n63) & (!n979)) + ((!n23) & (!n64) & (n63) & (n979)) + ((!n23) & (n64) & (!n63) & (n979)) + ((!n23) & (n64) & (n63) & (!n979)) + ((!n23) & (n64) & (n63) & (n979)) + ((n23) & (n64) & (!n63) & (n979)) + ((n23) & (n64) & (n63) & (!n979)) + ((n23) & (n64) & (n63) & (n979)));
	assign n1050 = (((!i_19_) & (!n163) & (!n347)) + ((!i_19_) & (!n163) & (n347)) + ((!i_19_) & (n163) & (!n347)) + ((!i_19_) & (n163) & (n347)) + ((i_19_) & (!n163) & (n347)) + ((i_19_) & (n163) & (!n347)) + ((i_19_) & (n163) & (n347)));
	assign n1049 = (((n1050) & (!i_28_) & (!n345) & (n199)) + ((n1050) & (!i_28_) & (n345) & (!n199)) + ((n1050) & (!i_28_) & (n345) & (n199)) + ((n1050) & (i_28_) & (!n345) & (!n199)) + ((n1050) & (i_28_) & (!n345) & (n199)) + ((n1050) & (i_28_) & (n345) & (!n199)) + ((n1050) & (i_28_) & (n345) & (n199)));
	assign n1051 = (((!n195) & (n200) & (!n356) & (!n382)) + ((!n195) & (n200) & (n356) & (!n382)) + ((n195) & (!n200) & (!n356) & (!n382)) + ((n195) & (n200) & (!n356) & (!n382)) + ((n195) & (n200) & (n356) & (!n382)));
	assign n1053 = (((!n121) & (!n190) & (!n378) & (!n611)) + ((!n121) & (!n190) & (!n378) & (n611)) + ((!n121) & (n190) & (!n378) & (!n611)) + ((!n121) & (n190) & (!n378) & (n611)) + ((n121) & (!n190) & (!n378) & (n611)) + ((n121) & (n190) & (!n378) & (!n611)) + ((n121) & (n190) & (!n378) & (n611)));
	assign n1055 = (((!n11) & (!n86) & (!n375) & (n377)) + ((!n11) & (!n86) & (n375) & (n377)) + ((!n11) & (n86) & (!n375) & (!n377)) + ((!n11) & (n86) & (!n375) & (n377)) + ((!n11) & (n86) & (n375) & (!n377)) + ((!n11) & (n86) & (n375) & (n377)) + ((n11) & (!n86) & (n375) & (n377)) + ((n11) & (n86) & (n375) & (!n377)) + ((n11) & (n86) & (n375) & (n377)));
	assign n1057 = (((n1018) & (n63)));
	assign n1056 = (((!n143) & (!n168) & (!n356) & (n1057)) + ((!n143) & (n168) & (!n356) & (!n1057)) + ((!n143) & (n168) & (!n356) & (n1057)) + ((n143) & (!n168) & (!n356) & (n1057)) + ((n143) & (!n168) & (n356) & (n1057)) + ((n143) & (n168) & (!n356) & (!n1057)) + ((n143) & (n168) & (!n356) & (n1057)) + ((n143) & (n168) & (n356) & (!n1057)) + ((n143) & (n168) & (n356) & (n1057)));
	assign n1058 = (((!n78) & (n344) & (!n385) & (n1056)) + ((n78) & (!n344) & (!n385) & (n1056)) + ((n78) & (n344) & (!n385) & (n1056)));
	assign n1060 = (((!n95) & (!n331) & (n841)) + ((!n95) & (n331) & (n841)) + ((n95) & (n331) & (n841)));
	assign n1062 = (((!n130) & (!n304) & (n963) & (!n978)) + ((!n130) & (!n304) & (n963) & (n978)) + ((!n130) & (n304) & (n963) & (n978)) + ((n130) & (!n304) & (!n963) & (!n978)) + ((n130) & (!n304) & (!n963) & (n978)) + ((n130) & (!n304) & (n963) & (!n978)) + ((n130) & (!n304) & (n963) & (n978)) + ((n130) & (n304) & (!n963) & (n978)) + ((n130) & (n304) & (n963) & (n978)));
	assign n1063 = (((!n92) & (!n170) & (!n337) & (!n832)) + ((!n92) & (n170) & (!n337) & (!n832)) + ((!n92) & (n170) & (!n337) & (n832)) + ((n92) & (!n170) & (!n337) & (!n832)) + ((n92) & (!n170) & (!n337) & (n832)) + ((n92) & (n170) & (!n337) & (!n832)) + ((n92) & (n170) & (!n337) & (n832)));
	assign n1065 = (((!n91) & (n130)) + ((n91) & (!n130)) + ((n91) & (n130)));
	assign n1066 = (((!n121) & (!n241) & (!n304) & (!n648)) + ((!n121) & (!n241) & (!n304) & (n648)) + ((!n121) & (!n241) & (n304) & (n648)) + ((!n121) & (n241) & (!n304) & (!n648)) + ((!n121) & (n241) & (!n304) & (n648)) + ((!n121) & (n241) & (n304) & (n648)) + ((n121) & (n241) & (!n304) & (!n648)) + ((n121) & (n241) & (!n304) & (n648)) + ((n121) & (n241) & (n304) & (n648)));
	assign n1068 = (((!i_28_) & (!n229) & (!n611)) + ((!i_28_) & (!n229) & (n611)) + ((!i_28_) & (n229) & (n611)) + ((i_28_) & (!n229) & (!n611)) + ((i_28_) & (!n229) & (n611)) + ((i_28_) & (n229) & (!n611)) + ((i_28_) & (n229) & (n611)));
	assign n1067 = (((!i_7_) & (!n350) & (!n968) & (n1068)) + ((!i_7_) & (!n350) & (n968) & (n1068)) + ((!i_7_) & (n350) & (n968) & (n1068)) + ((i_7_) & (!n350) & (!n968) & (n1068)) + ((i_7_) & (!n350) & (n968) & (n1068)) + ((i_7_) & (n350) & (!n968) & (n1068)) + ((i_7_) & (n350) & (n968) & (n1068)));
	assign n1070 = (((!n313) & (n347)));
	assign n1069 = (((!n1070) & (n283) & (!n65) & (n240)) + ((!n1070) & (n283) & (n65) & (!n240)) + ((!n1070) & (n283) & (n65) & (n240)) + ((n1070) & (!n283) & (!n65) & (n240)) + ((n1070) & (!n283) & (n65) & (!n240)) + ((n1070) & (!n283) & (n65) & (n240)) + ((n1070) & (n283) & (!n65) & (n240)) + ((n1070) & (n283) & (n65) & (!n240)) + ((n1070) & (n283) & (n65) & (n240)));
	assign n1072 = (((!n170) & (!n101) & (!n92) & (n163)) + ((!n170) & (!n101) & (n92) & (!n163)) + ((!n170) & (!n101) & (n92) & (n163)) + ((!n170) & (n101) & (!n92) & (!n163)) + ((!n170) & (n101) & (!n92) & (n163)) + ((!n170) & (n101) & (n92) & (!n163)) + ((!n170) & (n101) & (n92) & (n163)) + ((n170) & (!n101) & (!n92) & (!n163)) + ((n170) & (!n101) & (!n92) & (n163)) + ((n170) & (!n101) & (n92) & (!n163)) + ((n170) & (!n101) & (n92) & (n163)) + ((n170) & (n101) & (!n92) & (!n163)) + ((n170) & (n101) & (!n92) & (n163)) + ((n170) & (n101) & (n92) & (!n163)) + ((n170) & (n101) & (n92) & (n163)));
	assign n1071 = (((!i_25_) & (!i_28_) & (!n1060) & (n1072)) + ((!i_25_) & (i_28_) & (!n1060) & (n1072)) + ((!i_25_) & (i_28_) & (n1060) & (n1072)) + ((i_25_) & (!i_28_) & (!n1060) & (n1072)) + ((i_25_) & (!i_28_) & (n1060) & (n1072)) + ((i_25_) & (i_28_) & (!n1060) & (n1072)) + ((i_25_) & (i_28_) & (n1060) & (n1072)));
	assign n1073 = (((!i_35_) & (!n69) & (!n339) & (n1071)) + ((!i_35_) & (!n69) & (n339) & (n1071)) + ((!i_35_) & (n69) & (!n339) & (n1071)) + ((!i_35_) & (n69) & (n339) & (n1071)) + ((i_35_) & (!n69) & (n339) & (n1071)) + ((i_35_) & (n69) & (!n339) & (n1071)) + ((i_35_) & (n69) & (n339) & (n1071)));
	assign n1074 = (((!n243) & (n342) & (!n348) & (n1073)) + ((n243) & (!n342) & (!n348) & (n1073)) + ((n243) & (n342) & (!n348) & (n1073)));
	assign n1076 = (((!n133) & (n249) & (!n352) & (!n355)) + ((n133) & (!n249) & (!n352) & (!n355)) + ((n133) & (n249) & (!n352) & (!n355)));
	assign n1079 = (((!n248) & (n332) & (!n358) & (n1076)) + ((n248) & (!n332) & (!n358) & (n1076)) + ((n248) & (n332) & (!n358) & (n1076)));
	assign n1082 = (((!i_30_) & (!n313) & (!n414)) + ((!i_30_) & (!n313) & (n414)) + ((!i_30_) & (n313) & (!n414)) + ((i_30_) & (!n313) & (!n414)) + ((i_30_) & (!n313) & (n414)) + ((i_30_) & (n313) & (!n414)) + ((i_30_) & (n313) & (n414)));
	assign n1081 = (((!n32) & (!n347) & (n1082)) + ((!n32) & (n347) & (n1082)) + ((n32) & (n347) & (n1082)));
	assign n1083 = (((!i_24_) & (!n26) & (!n367) & (n996)) + ((!i_24_) & (!n26) & (n367) & (n996)) + ((!i_24_) & (n26) & (!n367) & (n996)) + ((i_24_) & (!n26) & (!n367) & (!n996)) + ((i_24_) & (!n26) & (!n367) & (n996)) + ((i_24_) & (!n26) & (n367) & (!n996)) + ((i_24_) & (!n26) & (n367) & (n996)) + ((i_24_) & (n26) & (!n367) & (!n996)) + ((i_24_) & (n26) & (!n367) & (n996)));
	assign n1084 = (((!n11) & (!n283) & (!n308) & (!n414)) + ((!n11) & (!n283) & (!n308) & (n414)) + ((!n11) & (n283) & (!n308) & (!n414)) + ((!n11) & (n283) & (!n308) & (n414)) + ((!n11) & (n283) & (n308) & (!n414)) + ((!n11) & (n283) & (n308) & (n414)) + ((n11) & (!n283) & (!n308) & (!n414)) + ((n11) & (n283) & (!n308) & (!n414)) + ((n11) & (n283) & (n308) & (!n414)));
	assign n1085 = (((!n317) & (!n322) & (!n1083) & (!n1084)) + ((!n317) & (!n322) & (!n1083) & (n1084)) + ((!n317) & (!n322) & (n1083) & (!n1084)) + ((!n317) & (!n322) & (n1083) & (n1084)) + ((!n317) & (n322) & (n1083) & (n1084)));
	assign n1087 = (((!i_13_) & (i_24_)) + ((i_13_) & (!i_24_)) + ((i_13_) & (i_24_)));
	assign n1088 = (((!n191) & (n1087) & (!n194) & (n145)) + ((!n191) & (n1087) & (n194) & (!n145)) + ((!n191) & (n1087) & (n194) & (n145)) + ((n191) & (!n1087) & (!n194) & (n145)) + ((n191) & (!n1087) & (n194) & (!n145)) + ((n191) & (!n1087) & (n194) & (n145)) + ((n191) & (n1087) & (!n194) & (n145)) + ((n191) & (n1087) & (n194) & (!n145)) + ((n191) & (n1087) & (n194) & (n145)));
	assign n1089 = (((!n127) & (!n256) & (!n274) & (!n997)) + ((!n127) & (!n256) & (!n274) & (n997)) + ((!n127) & (n256) & (!n274) & (n997)) + ((n127) & (!n256) & (!n274) & (!n997)) + ((n127) & (!n256) & (!n274) & (n997)) + ((n127) & (n256) & (!n274) & (!n997)) + ((n127) & (n256) & (!n274) & (n997)));
	assign n1092 = (((!i_2_) & (!n22) & (!n49)) + ((!i_2_) & (!n22) & (n49)) + ((!i_2_) & (n22) & (n49)) + ((i_2_) & (!n22) & (!n49)) + ((i_2_) & (!n22) & (n49)) + ((i_2_) & (n22) & (!n49)) + ((i_2_) & (n22) & (n49)));
	assign n1091 = (((n1092) & (!i_13_) & (!i_3_) & (n198)) + ((n1092) & (!i_13_) & (i_3_) & (!n198)) + ((n1092) & (!i_13_) & (i_3_) & (n198)) + ((n1092) & (i_13_) & (!i_3_) & (!n198)) + ((n1092) & (i_13_) & (!i_3_) & (n198)) + ((n1092) & (i_13_) & (i_3_) & (!n198)) + ((n1092) & (i_13_) & (i_3_) & (n198)));
	assign n1094 = (((!n136) & (!n189) & (!n229)) + ((!n136) & (n189) & (!n229)) + ((!n136) & (n189) & (n229)) + ((n136) & (!n189) & (!n229)) + ((n136) & (!n189) & (n229)) + ((n136) & (n189) & (!n229)) + ((n136) & (n189) & (n229)));
	assign n1093 = (((!i_12_) & (!n273) & (!n278) & (n1094)) + ((!i_12_) & (n273) & (!n278) & (n1094)) + ((i_12_) & (n273) & (!n278) & (n1094)));
	assign n1097 = (((!i_26_) & (!n35) & (!n841) & (!n1002)) + ((!i_26_) & (!n35) & (!n841) & (n1002)) + ((!i_26_) & (!n35) & (n841) & (!n1002)) + ((i_26_) & (!n35) & (!n841) & (!n1002)) + ((i_26_) & (!n35) & (!n841) & (n1002)) + ((i_26_) & (!n35) & (n841) & (!n1002)) + ((i_26_) & (n35) & (!n841) & (!n1002)) + ((i_26_) & (n35) & (!n841) & (n1002)) + ((i_26_) & (n35) & (n841) & (!n1002)));
	assign n1100 = (((!n146) & (!n240) & (n162)) + ((!n146) & (n240) & (!n162)) + ((!n146) & (n240) & (n162)) + ((n146) & (!n240) & (!n162)) + ((n146) & (!n240) & (n162)) + ((n146) & (n240) & (!n162)) + ((n146) & (n240) & (n162)));
	assign n1099 = (((n1100) & (!i_28_) & (!n242) & (n124)) + ((n1100) & (!i_28_) & (n242) & (!n124)) + ((n1100) & (!i_28_) & (n242) & (n124)) + ((n1100) & (i_28_) & (!n242) & (!n124)) + ((n1100) & (i_28_) & (!n242) & (n124)) + ((n1100) & (i_28_) & (n242) & (!n124)) + ((n1100) & (i_28_) & (n242) & (n124)));
	assign n1101 = (((!i_23_) & (!n237) & (!n356) & (n957)) + ((!i_23_) & (!n237) & (n356) & (n957)) + ((!i_23_) & (n237) & (!n356) & (!n957)) + ((!i_23_) & (n237) & (!n356) & (n957)) + ((!i_23_) & (n237) & (n356) & (!n957)) + ((!i_23_) & (n237) & (n356) & (n957)) + ((i_23_) & (!n237) & (!n356) & (n957)) + ((i_23_) & (n237) & (!n356) & (!n957)) + ((i_23_) & (n237) & (!n356) & (n957)));
	assign n1102 = (((!n53) & (!n230) & (!n282) & (!n279)) + ((!n53) & (!n230) & (!n282) & (n279)) + ((!n53) & (!n230) & (n282) & (!n279)) + ((n53) & (!n230) & (!n282) & (!n279)) + ((n53) & (!n230) & (!n282) & (n279)) + ((n53) & (!n230) & (n282) & (!n279)) + ((n53) & (!n230) & (n282) & (n279)));
	assign n1107 = (((!i_18_) & (!i_24_) & (!n191)) + ((!i_18_) & (!i_24_) & (n191)) + ((!i_18_) & (i_24_) & (!n191)) + ((!i_18_) & (i_24_) & (n191)) + ((i_18_) & (!i_24_) & (n191)) + ((i_18_) & (i_24_) & (!n191)) + ((i_18_) & (i_24_) & (n191)));
	assign n1106 = (((n1107) & (!n194) & (n144)) + ((n1107) & (n194) & (!n144)) + ((n1107) & (n194) & (n144)));
	assign n1108 = (((!n163) & (!n207) & (!n350) & (n995)) + ((!n163) & (n207) & (!n350) & (n995)) + ((!n163) & (n207) & (n350) & (n995)) + ((n163) & (!n207) & (!n350) & (!n995)) + ((n163) & (!n207) & (!n350) & (n995)) + ((n163) & (n207) & (!n350) & (!n995)) + ((n163) & (n207) & (!n350) & (n995)) + ((n163) & (n207) & (n350) & (!n995)) + ((n163) & (n207) & (n350) & (n995)));
	assign n1109 = (((!i_9_) & (!n36) & (!n41) & (!n45)) + ((!i_9_) & (n36) & (!n41) & (!n45)) + ((i_9_) & (n36) & (!n41) & (!n45)));
	assign n1112 = (((!n39) & (n147) & (!n256) & (!n1000)) + ((!n39) & (n147) & (!n256) & (n1000)) + ((!n39) & (n147) & (n256) & (n1000)) + ((n39) & (!n147) & (!n256) & (!n1000)) + ((n39) & (!n147) & (!n256) & (n1000)) + ((n39) & (!n147) & (n256) & (n1000)) + ((n39) & (n147) & (!n256) & (!n1000)) + ((n39) & (n147) & (!n256) & (n1000)) + ((n39) & (n147) & (n256) & (n1000)));
	assign n1114 = (((n1020) & (n454)));
	assign n1113 = (((!n1114) & (n173) & (!n69) & (n164)) + ((!n1114) & (n173) & (n69) & (!n164)) + ((!n1114) & (n173) & (n69) & (n164)) + ((n1114) & (!n173) & (!n69) & (n164)) + ((n1114) & (!n173) & (n69) & (!n164)) + ((n1114) & (!n173) & (n69) & (n164)) + ((n1114) & (n173) & (!n69) & (n164)) + ((n1114) & (n173) & (n69) & (!n164)) + ((n1114) & (n173) & (n69) & (n164)));
	assign n1115 = (((!n140) & (!n143) & (!n394) & (!n402)) + ((!n140) & (n143) & (!n394) & (!n402)) + ((!n140) & (n143) & (n394) & (!n402)) + ((n140) & (!n143) & (!n394) & (!n402)) + ((n140) & (!n143) & (!n394) & (n402)) + ((n140) & (n143) & (!n394) & (!n402)) + ((n140) & (n143) & (!n394) & (n402)) + ((n140) & (n143) & (n394) & (!n402)) + ((n140) & (n143) & (n394) & (n402)));
	assign n1116 = (((!i_31_) & (!n1127) & (n90)) + ((!i_31_) & (n1127) & (!n90)) + ((!i_31_) & (n1127) & (n90)) + ((i_31_) & (!n1127) & (!n90)) + ((i_31_) & (!n1127) & (n90)) + ((i_31_) & (n1127) & (!n90)) + ((i_31_) & (n1127) & (n90)));
	assign n1117 = (((!i_2_) & (!i_8_) & (!n135) & (!n394)) + ((!i_2_) & (!i_8_) & (n135) & (!n394)) + ((!i_2_) & (!i_8_) & (n135) & (n394)) + ((!i_2_) & (i_8_) & (!n135) & (!n394)) + ((!i_2_) & (i_8_) & (!n135) & (n394)) + ((!i_2_) & (i_8_) & (n135) & (!n394)) + ((!i_2_) & (i_8_) & (n135) & (n394)) + ((i_2_) & (!i_8_) & (!n135) & (!n394)) + ((i_2_) & (!i_8_) & (!n135) & (n394)) + ((i_2_) & (!i_8_) & (n135) & (!n394)) + ((i_2_) & (!i_8_) & (n135) & (n394)) + ((i_2_) & (i_8_) & (!n135) & (!n394)) + ((i_2_) & (i_8_) & (!n135) & (n394)) + ((i_2_) & (i_8_) & (n135) & (!n394)) + ((i_2_) & (i_8_) & (n135) & (n394)));
	assign n1120 = (((!i_34_) & (!n531) & (!n680)) + ((!i_34_) & (!n531) & (n680)) + ((!i_34_) & (n531) & (!n680)) + ((!i_34_) & (n531) & (n680)) + ((i_34_) & (!n531) & (!n680)) + ((i_34_) & (!n531) & (n680)) + ((i_34_) & (n531) & (n680)));
	assign n1118 = (((!n78) & (!n107) & (!n394) & (n1120)) + ((!n78) & (!n107) & (n394) & (n1120)) + ((!n78) & (n107) & (!n394) & (n1120)) + ((n78) & (!n107) & (!n394) & (n1120)) + ((n78) & (!n107) & (n394) & (n1120)) + ((n78) & (n107) & (!n394) & (n1120)) + ((n78) & (n107) & (n394) & (n1120)));
	assign n1122 = (((!n89) & (!n97) & (n148)) + ((!n89) & (n97) & (!n148)) + ((!n89) & (n97) & (n148)) + ((n89) & (!n97) & (!n148)) + ((n89) & (!n97) & (n148)) + ((n89) & (n97) & (!n148)) + ((n89) & (n97) & (n148)));
	assign n1121 = (((!i_13_) & (!n85) & (!n371) & (n1122)) + ((!i_13_) & (!n85) & (n371) & (n1122)) + ((!i_13_) & (n85) & (!n371) & (n1122)) + ((!i_13_) & (n85) & (n371) & (n1122)) + ((i_13_) & (!n85) & (n371) & (n1122)) + ((i_13_) & (n85) & (!n371) & (n1122)) + ((i_13_) & (n85) & (n371) & (n1122)));
	assign n1124 = (((!i_2_) & (!n972) & (n131)) + ((!i_2_) & (n972) & (!n131)) + ((!i_2_) & (n972) & (n131)) + ((i_2_) & (!n972) & (!n131)) + ((i_2_) & (!n972) & (n131)) + ((i_2_) & (n972) & (!n131)) + ((i_2_) & (n972) & (n131)));
	assign n1123 = (((!n86) & (n102) & (!n105) & (n1124)) + ((n86) & (!n102) & (!n105) & (n1124)) + ((n86) & (n102) & (!n105) & (n1124)));
	assign n1128 = (((!i_2_) & (!i_8_) & (!i_31_) & (!n306)) + ((!i_2_) & (!i_8_) & (i_31_) & (!n306)) + ((!i_2_) & (!i_8_) & (i_31_) & (n306)) + ((!i_2_) & (i_8_) & (!i_31_) & (!n306)) + ((!i_2_) & (i_8_) & (!i_31_) & (n306)) + ((!i_2_) & (i_8_) & (i_31_) & (!n306)) + ((!i_2_) & (i_8_) & (i_31_) & (n306)) + ((i_2_) & (!i_8_) & (!i_31_) & (!n306)) + ((i_2_) & (!i_8_) & (!i_31_) & (n306)) + ((i_2_) & (!i_8_) & (i_31_) & (!n306)) + ((i_2_) & (!i_8_) & (i_31_) & (n306)) + ((i_2_) & (i_8_) & (!i_31_) & (!n306)) + ((i_2_) & (i_8_) & (!i_31_) & (n306)) + ((i_2_) & (i_8_) & (i_31_) & (!n306)) + ((i_2_) & (i_8_) & (i_31_) & (n306)));
	assign n1127 = (((n1014) & (n40)));
	assign n1126 = (((!n394) & (!n972) & (n1128) & (!n1127)) + ((!n394) & (!n972) & (n1128) & (n1127)) + ((!n394) & (n972) & (n1128) & (!n1127)) + ((!n394) & (n972) & (n1128) & (n1127)) + ((n394) & (!n972) & (n1128) & (n1127)) + ((n394) & (n972) & (n1128) & (!n1127)) + ((n394) & (n972) & (n1128) & (n1127)));
	assign n1130 = (((!i_10_) & (!n61) & (!n402)) + ((!i_10_) & (n61) & (!n402)) + ((!i_10_) & (n61) & (n402)) + ((i_10_) & (!n61) & (!n402)) + ((i_10_) & (!n61) & (n402)) + ((i_10_) & (n61) & (!n402)) + ((i_10_) & (n61) & (n402)));
	assign n1129 = (((!i_29_) & (!n1002) & (!n1003) & (n1130)) + ((!i_29_) & (!n1002) & (n1003) & (n1130)) + ((!i_29_) & (n1002) & (!n1003) & (n1130)) + ((!i_29_) & (n1002) & (n1003) & (n1130)) + ((i_29_) & (!n1002) & (n1003) & (n1130)));
	assign n1131 = (((!n968) & (n1001) & (!n57) & (n326)) + ((!n968) & (n1001) & (n57) & (!n326)) + ((!n968) & (n1001) & (n57) & (n326)) + ((n968) & (!n1001) & (!n57) & (n326)) + ((n968) & (!n1001) & (n57) & (!n326)) + ((n968) & (!n1001) & (n57) & (n326)) + ((n968) & (n1001) & (!n57) & (n326)) + ((n968) & (n1001) & (n57) & (!n326)) + ((n968) & (n1001) & (n57) & (n326)));
	assign n1132 = (((!n68) & (!n322) & (n1131)) + ((n68) & (!n322) & (n1131)) + ((n68) & (n322) & (n1131)));
	assign n1134 = (((!n253) & (!n531) & (!n680)) + ((!n253) & (!n531) & (n680)) + ((!n253) & (n531) & (!n680)) + ((!n253) & (n531) & (n680)) + ((n253) & (!n531) & (!n680)) + ((n253) & (!n531) & (n680)) + ((n253) & (n531) & (n680)));
	assign n1133 = (((!n44) & (!n49) & (!n969) & (n1134)) + ((!n44) & (!n49) & (n969) & (n1134)) + ((!n44) & (n49) & (!n969) & (n1134)) + ((!n44) & (n49) & (n969) & (n1134)) + ((n44) & (!n49) & (n969) & (n1134)) + ((n44) & (n49) & (!n969) & (n1134)) + ((n44) & (n49) & (n969) & (n1134)));
	assign n1135 = (((!i_9_) & (!i_12_) & (!n53) & (n1133)) + ((!i_9_) & (!i_12_) & (n53) & (n1133)) + ((!i_9_) & (i_12_) & (!n53) & (n1133)) + ((!i_9_) & (i_12_) & (n53) & (n1133)) + ((i_9_) & (!i_12_) & (!n53) & (n1133)) + ((i_9_) & (!i_12_) & (n53) & (n1133)) + ((i_9_) & (i_12_) & (n53) & (n1133)));
	assign n1136 = (((!n109) & (!n113) & (!n117) & (!n324)) + ((n109) & (!n113) & (!n117) & (!n324)) + ((n109) & (!n113) & (!n117) & (n324)));
	assign n1140 = (((!n89) & (!n147) & (!n429)) + ((!n89) & (n147) & (!n429)) + ((!n89) & (n147) & (n429)) + ((n89) & (!n147) & (!n429)) + ((n89) & (!n147) & (n429)) + ((n89) & (n147) & (!n429)) + ((n89) & (n147) & (n429)));
	assign n1139 = (((n1140) & (!n140) & (!n1070) & (n162)) + ((n1140) & (!n140) & (n1070) & (!n162)) + ((n1140) & (!n140) & (n1070) & (n162)) + ((n1140) & (n140) & (!n1070) & (!n162)) + ((n1140) & (n140) & (!n1070) & (n162)) + ((n1140) & (n140) & (n1070) & (!n162)) + ((n1140) & (n140) & (n1070) & (n162)));
	assign n1141 = (((!i_35_) & (!n186) & (n139)) + ((!i_35_) & (n186) & (!n139)) + ((!i_35_) & (n186) & (n139)) + ((i_35_) & (!n186) & (!n139)) + ((i_35_) & (!n186) & (n139)) + ((i_35_) & (n186) & (!n139)) + ((i_35_) & (n186) & (n139)));
	assign n1143 = (((!i_38_) & (!n403) & (!n1074) & (!n1079)) + ((!i_38_) & (!n403) & (!n1074) & (n1079)) + ((!i_38_) & (!n403) & (n1074) & (!n1079)) + ((!i_38_) & (!n403) & (n1074) & (n1079)) + ((i_38_) & (!n403) & (n1074) & (n1079)));
	assign n1147 = (((n300) & (!n301) & (!n305) & (!n309) & (n314) & (n1085) & (n1226) & (n1264)));
	assign n1146 = (((!i_29_) & (!i_34_) & (n319) & (!n1147)) + ((!i_29_) & (!i_34_) & (n319) & (n1147)) + ((!i_29_) & (i_34_) & (n319) & (n1147)) + ((i_29_) & (!i_34_) & (!n319) & (!n1147)) + ((i_29_) & (!i_34_) & (!n319) & (n1147)) + ((i_29_) & (!i_34_) & (n319) & (!n1147)) + ((i_29_) & (!i_34_) & (n319) & (n1147)) + ((i_29_) & (i_34_) & (!n319) & (n1147)) + ((i_29_) & (i_34_) & (n319) & (n1147)));
	assign n1149 = (((!n10) & (!n408) & (!n412) & (!n998)) + ((!n10) & (!n408) & (!n412) & (n998)) + ((n10) & (!n408) & (!n412) & (n998)));
	assign n1152 = (((!n127) & (n264) & (!n122) & (n260)) + ((!n127) & (n264) & (n122) & (!n260)) + ((!n127) & (n264) & (n122) & (n260)) + ((n127) & (!n264) & (!n122) & (n260)) + ((n127) & (!n264) & (n122) & (!n260)) + ((n127) & (!n264) & (n122) & (n260)) + ((n127) & (n264) & (!n122) & (n260)) + ((n127) & (n264) & (n122) & (!n260)) + ((n127) & (n264) & (n122) & (n260)));
	assign n1153 = (((!i_24_) & (!n415) & (n1099) & (n1101)) + ((i_24_) & (!n415) & (!n1099) & (!n1101)) + ((i_24_) & (!n415) & (!n1099) & (n1101)) + ((i_24_) & (!n415) & (n1099) & (!n1101)) + ((i_24_) & (!n415) & (n1099) & (n1101)));
	assign n1155 = (((!n205) & (!n425) & (n1109) & (n1112)) + ((n205) & (!n425) & (!n1109) & (!n1112)) + ((n205) & (!n425) & (!n1109) & (n1112)) + ((n205) & (!n425) & (n1109) & (!n1112)) + ((n205) & (!n425) & (n1109) & (n1112)));
	assign n1157 = (((!n198) & (!n428) & (n979) & (n1155)) + ((n198) & (!n428) & (!n979) & (n1155)) + ((n198) & (!n428) & (n979) & (n1155)));
	assign n1159 = (((!n157) & (n195) & (!n132) & (n265)) + ((!n157) & (n195) & (n132) & (!n265)) + ((!n157) & (n195) & (n132) & (n265)) + ((n157) & (!n195) & (!n132) & (n265)) + ((n157) & (!n195) & (n132) & (!n265)) + ((n157) & (!n195) & (n132) & (n265)) + ((n157) & (n195) & (!n132) & (n265)) + ((n157) & (n195) & (n132) & (!n265)) + ((n157) & (n195) & (n132) & (n265)));
	assign n1160 = (((n217) & (!i_22_) & (n1136) & (n1135)) + ((n217) & (i_22_) & (!n1136) & (!n1135)) + ((n217) & (i_22_) & (!n1136) & (n1135)) + ((n217) & (i_22_) & (n1136) & (!n1135)) + ((n217) & (i_22_) & (n1136) & (n1135)));
	assign n1163 = (((!n1012) & (n558)) + ((n1012) & (!n558)) + ((n1012) & (n558)));
	assign n1164 = (((!n59) & (!n447) & (!n481) & (!n1261)) + ((!n59) & (!n447) & (!n481) & (n1261)) + ((!n59) & (!n447) & (n481) & (!n1261)) + ((n59) & (!n447) & (!n481) & (!n1261)) + ((n59) & (!n447) & (n481) & (!n1261)));
	assign n1169 = (((!n1018) & (n1019)) + ((n1018) & (!n1019)) + ((n1018) & (n1019)));
	assign n1171 = (((!n213) & (!n253) & (!n315)) + ((!n213) & (!n253) & (n315)) + ((!n213) & (n253) & (n315)) + ((n213) & (!n253) & (!n315)) + ((n213) & (!n253) & (n315)) + ((n213) & (n253) & (!n315)) + ((n213) & (n253) & (n315)));
	assign n1170 = (((!i_20_) & (!n722) & (!n1003) & (n1171)) + ((!i_20_) & (!n722) & (n1003) & (n1171)) + ((!i_20_) & (n722) & (!n1003) & (n1171)) + ((!i_20_) & (n722) & (n1003) & (n1171)) + ((i_20_) & (!n722) & (!n1003) & (n1171)) + ((i_20_) & (n722) & (!n1003) & (n1171)) + ((i_20_) & (n722) & (n1003) & (n1171)));
	assign n1173 = (((!i_31_) & (!n715) & (!n974)) + ((!i_31_) & (!n715) & (n974)) + ((!i_31_) & (n715) & (!n974)) + ((!i_31_) & (n715) & (n974)) + ((i_31_) & (!n715) & (n974)) + ((i_31_) & (n715) & (!n974)) + ((i_31_) & (n715) & (n974)));
	assign n1172 = (((n1173) & (!n642) & (!n340) & (n717)) + ((n1173) & (!n642) & (n340) & (!n717)) + ((n1173) & (!n642) & (n340) & (n717)) + ((n1173) & (n642) & (!n340) & (!n717)) + ((n1173) & (n642) & (!n340) & (n717)) + ((n1173) & (n642) & (n340) & (!n717)) + ((n1173) & (n642) & (n340) & (n717)));
	assign n1174 = (((!i_7_) & (!n972) & (n993)) + ((!i_7_) & (n972) & (!n993)) + ((!i_7_) & (n972) & (n993)) + ((i_7_) & (!n972) & (!n993)) + ((i_7_) & (!n972) & (n993)) + ((i_7_) & (n972) & (!n993)) + ((i_7_) & (n972) & (n993)));
	assign n1175 = (((!n245) & (!n667) & (!n1025) & (!n1026)) + ((!n245) & (!n667) & (!n1025) & (n1026)) + ((!n245) & (!n667) & (n1025) & (!n1026)) + ((!n245) & (!n667) & (n1025) & (n1026)) + ((n245) & (!n667) & (!n1025) & (n1026)) + ((n245) & (!n667) & (n1025) & (!n1026)) + ((n245) & (!n667) & (n1025) & (n1026)));
	assign n1179 = (((!n1012) & (n1019)) + ((n1012) & (!n1019)) + ((n1012) & (n1019)));
	assign n1180 = (((!n649) & (!n1028) & (!n345) & (n556)) + ((!n649) & (!n1028) & (n345) & (!n556)) + ((!n649) & (!n1028) & (n345) & (n556)) + ((!n649) & (n1028) & (!n345) & (!n556)) + ((!n649) & (n1028) & (!n345) & (n556)) + ((!n649) & (n1028) & (n345) & (!n556)) + ((!n649) & (n1028) & (n345) & (n556)) + ((n649) & (!n1028) & (!n345) & (!n556)) + ((n649) & (!n1028) & (!n345) & (n556)) + ((n649) & (!n1028) & (n345) & (!n556)) + ((n649) & (!n1028) & (n345) & (n556)) + ((n649) & (n1028) & (!n345) & (!n556)) + ((n649) & (n1028) & (!n345) & (n556)) + ((n649) & (n1028) & (n345) & (!n556)) + ((n649) & (n1028) & (n345) & (n556)));
	assign n1181 = (((!i_0_) & (!i_30_) & (!n229) & (!n477) & (!n664) & (!n1027)) + ((!i_0_) & (!i_30_) & (!n229) & (!n477) & (!n664) & (n1027)) + ((!i_0_) & (!i_30_) & (!n229) & (!n477) & (n664) & (!n1027)) + ((!i_0_) & (!i_30_) & (!n229) & (!n477) & (n664) & (n1027)) + ((!i_0_) & (!i_30_) & (!n229) & (n477) & (!n664) & (!n1027)) + ((!i_0_) & (!i_30_) & (!n229) & (n477) & (!n664) & (n1027)) + ((!i_0_) & (!i_30_) & (!n229) & (n477) & (n664) & (!n1027)) + ((!i_0_) & (!i_30_) & (!n229) & (n477) & (n664) & (n1027)) + ((!i_0_) & (!i_30_) & (n229) & (!n477) & (!n664) & (n1027)) + ((!i_0_) & (!i_30_) & (n229) & (!n477) & (n664) & (!n1027)) + ((!i_0_) & (!i_30_) & (n229) & (!n477) & (n664) & (n1027)) + ((!i_0_) & (!i_30_) & (n229) & (n477) & (!n664) & (!n1027)) + ((!i_0_) & (!i_30_) & (n229) & (n477) & (!n664) & (n1027)) + ((!i_0_) & (!i_30_) & (n229) & (n477) & (n664) & (!n1027)) + ((!i_0_) & (!i_30_) & (n229) & (n477) & (n664) & (n1027)) + ((!i_0_) & (i_30_) & (!n229) & (!n477) & (!n664) & (!n1027)) + ((!i_0_) & (i_30_) & (!n229) & (!n477) & (!n664) & (n1027)) + ((!i_0_) & (i_30_) & (!n229) & (!n477) & (n664) & (!n1027)) + ((!i_0_) & (i_30_) & (!n229) & (!n477) & (n664) & (n1027)) + ((!i_0_) & (i_30_) & (!n229) & (n477) & (!n664) & (!n1027)) + ((!i_0_) & (i_30_) & (!n229) & (n477) & (!n664) & (n1027)) + ((!i_0_) & (i_30_) & (!n229) & (n477) & (n664) & (!n1027)) + ((!i_0_) & (i_30_) & (!n229) & (n477) & (n664) & (n1027)) + ((!i_0_) & (i_30_) & (n229) & (!n477) & (!n664) & (!n1027)) + ((!i_0_) & (i_30_) & (n229) & (!n477) & (!n664) & (n1027)) + ((!i_0_) & (i_30_) & (n229) & (!n477) & (n664) & (!n1027)) + ((!i_0_) & (i_30_) & (n229) & (!n477) & (n664) & (n1027)) + ((!i_0_) & (i_30_) & (n229) & (n477) & (!n664) & (!n1027)) + ((!i_0_) & (i_30_) & (n229) & (n477) & (!n664) & (n1027)) + ((!i_0_) & (i_30_) & (n229) & (n477) & (n664) & (!n1027)) + ((!i_0_) & (i_30_) & (n229) & (n477) & (n664) & (n1027)) + ((i_0_) & (!i_30_) & (!n229) & (!n477) & (!n664) & (!n1027)) + ((i_0_) & (!i_30_) & (!n229) & (!n477) & (!n664) & (n1027)) + ((i_0_) & (!i_30_) & (!n229) & (!n477) & (n664) & (!n1027)) + ((i_0_) & (!i_30_) & (!n229) & (!n477) & (n664) & (n1027)) + ((i_0_) & (!i_30_) & (!n229) & (n477) & (!n664) & (!n1027)) + ((i_0_) & (!i_30_) & (!n229) & (n477) & (!n664) & (n1027)) + ((i_0_) & (!i_30_) & (!n229) & (n477) & (n664) & (!n1027)) + ((i_0_) & (!i_30_) & (!n229) & (n477) & (n664) & (n1027)) + ((i_0_) & (!i_30_) & (n229) & (!n477) & (!n664) & (!n1027)) + ((i_0_) & (!i_30_) & (n229) & (!n477) & (!n664) & (n1027)) + ((i_0_) & (!i_30_) & (n229) & (!n477) & (n664) & (!n1027)) + ((i_0_) & (!i_30_) & (n229) & (!n477) & (n664) & (n1027)) + ((i_0_) & (!i_30_) & (n229) & (n477) & (!n664) & (!n1027)) + ((i_0_) & (!i_30_) & (n229) & (n477) & (!n664) & (n1027)) + ((i_0_) & (!i_30_) & (n229) & (n477) & (n664) & (!n1027)) + ((i_0_) & (!i_30_) & (n229) & (n477) & (n664) & (n1027)) + ((i_0_) & (i_30_) & (!n229) & (!n477) & (!n664) & (!n1027)) + ((i_0_) & (i_30_) & (!n229) & (!n477) & (!n664) & (n1027)) + ((i_0_) & (i_30_) & (!n229) & (!n477) & (n664) & (!n1027)) + ((i_0_) & (i_30_) & (!n229) & (!n477) & (n664) & (n1027)) + ((i_0_) & (i_30_) & (!n229) & (n477) & (!n664) & (!n1027)) + ((i_0_) & (i_30_) & (!n229) & (n477) & (!n664) & (n1027)) + ((i_0_) & (i_30_) & (!n229) & (n477) & (n664) & (!n1027)) + ((i_0_) & (i_30_) & (!n229) & (n477) & (n664) & (n1027)) + ((i_0_) & (i_30_) & (n229) & (!n477) & (!n664) & (!n1027)) + ((i_0_) & (i_30_) & (n229) & (!n477) & (!n664) & (n1027)) + ((i_0_) & (i_30_) & (n229) & (!n477) & (n664) & (!n1027)) + ((i_0_) & (i_30_) & (n229) & (!n477) & (n664) & (n1027)) + ((i_0_) & (i_30_) & (n229) & (n477) & (!n664) & (!n1027)) + ((i_0_) & (i_30_) & (n229) & (n477) & (!n664) & (n1027)) + ((i_0_) & (i_30_) & (n229) & (n477) & (n664) & (!n1027)) + ((i_0_) & (i_30_) & (n229) & (n477) & (n664) & (n1027)));
	assign n1183 = (((!n442) & (!n1019) & (n559)) + ((!n442) & (n1019) & (!n559)) + ((!n442) & (n1019) & (n559)) + ((n442) & (!n1019) & (!n559)) + ((n442) & (!n1019) & (n559)) + ((n442) & (n1019) & (!n559)) + ((n442) & (n1019) & (n559)));
	assign n1182 = (((n1183) & (!n447) & (n618)) + ((n1183) & (n447) & (!n618)) + ((n1183) & (n447) & (n618)));
	assign n1186 = (((!i_7_) & (!i_23_) & (!n290) & (!n308) & (!n443)) + ((!i_7_) & (!i_23_) & (!n290) & (!n308) & (n443)) + ((!i_7_) & (!i_23_) & (!n290) & (n308) & (!n443)) + ((!i_7_) & (!i_23_) & (!n290) & (n308) & (n443)) + ((!i_7_) & (!i_23_) & (n290) & (!n308) & (!n443)) + ((!i_7_) & (!i_23_) & (n290) & (!n308) & (n443)) + ((!i_7_) & (!i_23_) & (n290) & (n308) & (n443)) + ((!i_7_) & (i_23_) & (!n290) & (!n308) & (!n443)) + ((!i_7_) & (i_23_) & (!n290) & (!n308) & (n443)) + ((!i_7_) & (i_23_) & (!n290) & (n308) & (!n443)) + ((!i_7_) & (i_23_) & (!n290) & (n308) & (n443)) + ((!i_7_) & (i_23_) & (n290) & (!n308) & (!n443)) + ((!i_7_) & (i_23_) & (n290) & (!n308) & (n443)) + ((!i_7_) & (i_23_) & (n290) & (n308) & (!n443)) + ((!i_7_) & (i_23_) & (n290) & (n308) & (n443)) + ((i_7_) & (!i_23_) & (!n290) & (!n308) & (!n443)) + ((i_7_) & (!i_23_) & (!n290) & (!n308) & (n443)) + ((i_7_) & (!i_23_) & (!n290) & (n308) & (!n443)) + ((i_7_) & (!i_23_) & (!n290) & (n308) & (n443)) + ((i_7_) & (!i_23_) & (n290) & (!n308) & (!n443)) + ((i_7_) & (!i_23_) & (n290) & (!n308) & (n443)) + ((i_7_) & (!i_23_) & (n290) & (n308) & (!n443)) + ((i_7_) & (!i_23_) & (n290) & (n308) & (n443)) + ((i_7_) & (i_23_) & (!n290) & (!n308) & (!n443)) + ((i_7_) & (i_23_) & (!n290) & (!n308) & (n443)) + ((i_7_) & (i_23_) & (!n290) & (n308) & (!n443)) + ((i_7_) & (i_23_) & (!n290) & (n308) & (n443)) + ((i_7_) & (i_23_) & (n290) & (!n308) & (!n443)) + ((i_7_) & (i_23_) & (n290) & (!n308) & (n443)) + ((i_7_) & (i_23_) & (n290) & (n308) & (!n443)) + ((i_7_) & (i_23_) & (n290) & (n308) & (n443)));
	assign n1187 = (((!n501) & (!n543) & (n646) & (!n1022)) + ((!n501) & (!n543) & (n646) & (n1022)) + ((!n501) & (n543) & (n646) & (n1022)) + ((n501) & (!n543) & (!n646) & (!n1022)) + ((n501) & (!n543) & (!n646) & (n1022)) + ((n501) & (!n543) & (n646) & (!n1022)) + ((n501) & (!n543) & (n646) & (n1022)) + ((n501) & (n543) & (!n646) & (n1022)) + ((n501) & (n543) & (n646) & (n1022)));
	assign n1189 = (((!i_37_) & (!n349) & (!n556) & (!n1028)) + ((!i_37_) & (!n349) & (!n556) & (n1028)) + ((!i_37_) & (!n349) & (n556) & (!n1028)) + ((!i_37_) & (!n349) & (n556) & (n1028)) + ((!i_37_) & (n349) & (!n556) & (!n1028)) + ((!i_37_) & (n349) & (!n556) & (n1028)) + ((!i_37_) & (n349) & (n556) & (!n1028)) + ((!i_37_) & (n349) & (n556) & (n1028)) + ((i_37_) & (!n349) & (!n556) & (!n1028)) + ((i_37_) & (!n349) & (!n556) & (n1028)) + ((i_37_) & (!n349) & (n556) & (!n1028)) + ((i_37_) & (!n349) & (n556) & (n1028)) + ((i_37_) & (n349) & (!n556) & (n1028)) + ((i_37_) & (n349) & (n556) & (!n1028)) + ((i_37_) & (n349) & (n556) & (n1028)));
	assign n1188 = (((!n376) & (!n543) & (!n612) & (n1189)) + ((!n376) & (!n543) & (n612) & (n1189)) + ((!n376) & (n543) & (n612) & (n1189)) + ((n376) & (!n543) & (!n612) & (n1189)) + ((n376) & (!n543) & (n612) & (n1189)) + ((n376) & (n543) & (!n612) & (n1189)) + ((n376) & (n543) & (n612) & (n1189)));
	assign n1191 = (((!i_2_) & (!i_16_) & (!n31)) + ((!i_2_) & (!i_16_) & (n31)) + ((!i_2_) & (i_16_) & (!n31)) + ((!i_2_) & (i_16_) & (n31)) + ((i_2_) & (!i_16_) & (n31)) + ((i_2_) & (i_16_) & (!n31)) + ((i_2_) & (i_16_) & (n31)));
	assign n1190 = (((n1191) & (!n502) & (!n84) & (n1015)) + ((n1191) & (!n502) & (n84) & (!n1015)) + ((n1191) & (!n502) & (n84) & (n1015)) + ((n1191) & (n502) & (!n84) & (!n1015)) + ((n1191) & (n502) & (!n84) & (n1015)) + ((n1191) & (n502) & (n84) & (!n1015)) + ((n1191) & (n502) & (n84) & (n1015)));
	assign n1192 = (((!i_37_) & (!n81) & (!n513) & (!n520)) + ((!i_37_) & (!n81) & (!n513) & (n520)) + ((!i_37_) & (!n81) & (n513) & (!n520)) + ((!i_37_) & (!n81) & (n513) & (n520)) + ((!i_37_) & (n81) & (!n513) & (!n520)) + ((!i_37_) & (n81) & (!n513) & (n520)) + ((!i_37_) & (n81) & (n513) & (!n520)) + ((!i_37_) & (n81) & (n513) & (n520)) + ((i_37_) & (!n81) & (!n513) & (n520)) + ((i_37_) & (!n81) & (n513) & (!n520)) + ((i_37_) & (!n81) & (n513) & (n520)) + ((i_37_) & (n81) & (!n513) & (!n520)) + ((i_37_) & (n81) & (!n513) & (n520)) + ((i_37_) & (n81) & (n513) & (!n520)) + ((i_37_) & (n81) & (n513) & (n520)));
	assign n1193 = (((!n347) & (!n350) & (!n514) & (n703)) + ((!n347) & (!n350) & (n514) & (n703)) + ((!n347) & (n350) & (n514) & (n703)) + ((n347) & (!n350) & (!n514) & (!n703)) + ((n347) & (!n350) & (!n514) & (n703)) + ((n347) & (!n350) & (n514) & (!n703)) + ((n347) & (!n350) & (n514) & (n703)) + ((n347) & (n350) & (n514) & (!n703)) + ((n347) & (n350) & (n514) & (n703)));
	assign n1195 = (((!i_30_) & (!i_31_) & (!n362) & (!n479)) + ((!i_30_) & (!i_31_) & (!n362) & (n479)) + ((!i_30_) & (!i_31_) & (n362) & (!n479)) + ((!i_30_) & (!i_31_) & (n362) & (n479)) + ((!i_30_) & (i_31_) & (!n362) & (!n479)) + ((!i_30_) & (i_31_) & (!n362) & (n479)) + ((!i_30_) & (i_31_) & (n362) & (n479)) + ((i_30_) & (!i_31_) & (!n362) & (!n479)) + ((i_30_) & (!i_31_) & (!n362) & (n479)) + ((i_30_) & (!i_31_) & (n362) & (!n479)) + ((i_30_) & (!i_31_) & (n362) & (n479)) + ((i_30_) & (i_31_) & (!n362) & (!n479)) + ((i_30_) & (i_31_) & (!n362) & (n479)) + ((i_30_) & (i_31_) & (n362) & (!n479)) + ((i_30_) & (i_31_) & (n362) & (n479)));
	assign n1194 = (((n1195) & (!i_14_) & (!n631) & (n461)) + ((n1195) & (!i_14_) & (n631) & (!n461)) + ((n1195) & (!i_14_) & (n631) & (n461)) + ((n1195) & (i_14_) & (!n631) & (!n461)) + ((n1195) & (i_14_) & (!n631) & (n461)) + ((n1195) & (i_14_) & (n631) & (!n461)) + ((n1195) & (i_14_) & (n631) & (n461)));
	assign n1197 = (((!n373) & (!n474) & (!n622) & (!n631) & (!n681)) + ((!n373) & (!n474) & (!n622) & (n631) & (!n681)) + ((!n373) & (!n474) & (!n622) & (n631) & (n681)) + ((!n373) & (!n474) & (n622) & (!n631) & (!n681)) + ((!n373) & (!n474) & (n622) & (!n631) & (n681)) + ((!n373) & (!n474) & (n622) & (n631) & (!n681)) + ((!n373) & (!n474) & (n622) & (n631) & (n681)) + ((!n373) & (n474) & (!n622) & (!n631) & (!n681)) + ((!n373) & (n474) & (!n622) & (!n631) & (n681)) + ((!n373) & (n474) & (!n622) & (n631) & (!n681)) + ((!n373) & (n474) & (!n622) & (n631) & (n681)) + ((!n373) & (n474) & (n622) & (!n631) & (!n681)) + ((!n373) & (n474) & (n622) & (!n631) & (n681)) + ((!n373) & (n474) & (n622) & (n631) & (!n681)) + ((!n373) & (n474) & (n622) & (n631) & (n681)) + ((n373) & (!n474) & (!n622) & (!n631) & (!n681)) + ((n373) & (!n474) & (!n622) & (!n631) & (n681)) + ((n373) & (!n474) & (!n622) & (n631) & (!n681)) + ((n373) & (!n474) & (!n622) & (n631) & (n681)) + ((n373) & (!n474) & (n622) & (!n631) & (!n681)) + ((n373) & (!n474) & (n622) & (!n631) & (n681)) + ((n373) & (!n474) & (n622) & (n631) & (!n681)) + ((n373) & (!n474) & (n622) & (n631) & (n681)) + ((n373) & (n474) & (!n622) & (!n631) & (!n681)) + ((n373) & (n474) & (!n622) & (!n631) & (n681)) + ((n373) & (n474) & (!n622) & (n631) & (!n681)) + ((n373) & (n474) & (!n622) & (n631) & (n681)) + ((n373) & (n474) & (n622) & (!n631) & (!n681)) + ((n373) & (n474) & (n622) & (!n631) & (n681)) + ((n373) & (n474) & (n622) & (n631) & (!n681)) + ((n373) & (n474) & (n622) & (n631) & (n681)));
	assign n1196 = (((!n452) & (!n543) & (!n813) & (n1197)) + ((!n452) & (!n543) & (n813) & (n1197)) + ((!n452) & (n543) & (n813) & (n1197)) + ((n452) & (!n543) & (!n813) & (n1197)) + ((n452) & (!n543) & (n813) & (n1197)) + ((n452) & (n543) & (!n813) & (n1197)) + ((n452) & (n543) & (n813) & (n1197)));
	assign n1198 = (((!n645) & (!n347) & (n572)) + ((!n645) & (n347) & (!n572)) + ((!n645) & (n347) & (n572)) + ((n645) & (!n347) & (!n572)) + ((n645) & (!n347) & (n572)) + ((n645) & (n347) & (!n572)) + ((n645) & (n347) & (n572)));
	assign n1200 = (((!n692) & (!n880) & (!n973)) + ((!n692) & (!n880) & (n973)) + ((!n692) & (n880) & (!n973)) + ((!n692) & (n880) & (n973)) + ((n692) & (!n880) & (!n973)) + ((n692) & (!n880) & (n973)) + ((n692) & (n880) & (n973)));
	assign n1199 = (((n1200) & (!n442) & (!n556) & (n1017)) + ((n1200) & (!n442) & (n556) & (!n1017)) + ((n1200) & (!n442) & (n556) & (n1017)) + ((n1200) & (n442) & (!n556) & (!n1017)) + ((n1200) & (n442) & (!n556) & (n1017)) + ((n1200) & (n442) & (n556) & (!n1017)) + ((n1200) & (n442) & (n556) & (n1017)));
	assign n1201 = (((!i_13_) & (!n624) & (n631)) + ((!i_13_) & (n624) & (!n631)) + ((!i_13_) & (n624) & (n631)) + ((i_13_) & (!n624) & (!n631)) + ((i_13_) & (!n624) & (n631)) + ((i_13_) & (n624) & (!n631)) + ((i_13_) & (n624) & (n631)));
	assign n1202 = (((!i_7_) & (!n550) & (n719) & (!n733)) + ((!i_7_) & (!n550) & (n719) & (n733)) + ((!i_7_) & (n550) & (!n719) & (!n733)) + ((!i_7_) & (n550) & (!n719) & (n733)) + ((!i_7_) & (n550) & (n719) & (!n733)) + ((!i_7_) & (n550) & (n719) & (n733)) + ((i_7_) & (!n550) & (n719) & (n733)) + ((i_7_) & (n550) & (!n719) & (n733)) + ((i_7_) & (n550) & (n719) & (n733)));
	assign n1203 = (((!n241) & (!n446) & (n695)) + ((!n241) & (n446) & (!n695)) + ((!n241) & (n446) & (n695)) + ((n241) & (!n446) & (!n695)) + ((n241) & (!n446) & (n695)) + ((n241) & (n446) & (!n695)) + ((n241) & (n446) & (n695)));
	assign n1204 = (((!n215) & (!n543) & (!n709) & (n713)) + ((!n215) & (!n543) & (n709) & (n713)) + ((!n215) & (n543) & (n709) & (n713)) + ((n215) & (!n543) & (!n709) & (!n713)) + ((n215) & (!n543) & (!n709) & (n713)) + ((n215) & (!n543) & (n709) & (!n713)) + ((n215) & (!n543) & (n709) & (n713)) + ((n215) & (n543) & (n709) & (!n713)) + ((n215) & (n543) & (n709) & (n713)));
	assign n1205 = (((!n697) & (n443) & (!n874) & (n674)) + ((!n697) & (n443) & (n874) & (!n674)) + ((!n697) & (n443) & (n874) & (n674)) + ((n697) & (!n443) & (!n874) & (n674)) + ((n697) & (!n443) & (n874) & (!n674)) + ((n697) & (!n443) & (n874) & (n674)) + ((n697) & (n443) & (!n874) & (n674)) + ((n697) & (n443) & (n874) & (!n674)) + ((n697) & (n443) & (n874) & (n674)));
	assign n1206 = (((!i_37_) & (!n290) & (!n634) & (!n658)) + ((!i_37_) & (!n290) & (!n634) & (n658)) + ((!i_37_) & (!n290) & (n634) & (!n658)) + ((!i_37_) & (!n290) & (n634) & (n658)) + ((!i_37_) & (n290) & (n634) & (!n658)) + ((!i_37_) & (n290) & (n634) & (n658)) + ((i_37_) & (!n290) & (!n634) & (n658)) + ((i_37_) & (!n290) & (n634) & (n658)) + ((i_37_) & (n290) & (n634) & (n658)));
	assign n1207 = (((!n613) & (n664) & (!i_14_) & (n582)) + ((!n613) & (n664) & (i_14_) & (!n582)) + ((!n613) & (n664) & (i_14_) & (n582)) + ((n613) & (!n664) & (!i_14_) & (n582)) + ((n613) & (!n664) & (i_14_) & (!n582)) + ((n613) & (!n664) & (i_14_) & (n582)) + ((n613) & (n664) & (!i_14_) & (n582)) + ((n613) & (n664) & (i_14_) & (!n582)) + ((n613) & (n664) & (i_14_) & (n582)));
	assign n1209 = (((!n529) & (n533) & (!n535) & (!n540) & (n998) & (n1268)));
	assign n1208 = (((!n10) & (!n362) & (!n567) & (!n1209)) + ((!n10) & (!n362) & (!n567) & (n1209)) + ((!n10) & (!n362) & (n567) & (!n1209)) + ((!n10) & (!n362) & (n567) & (n1209)) + ((!n10) & (n362) & (n567) & (!n1209)) + ((!n10) & (n362) & (n567) & (n1209)) + ((n10) & (!n362) & (!n567) & (n1209)) + ((n10) & (!n362) & (n567) & (n1209)) + ((n10) & (n362) & (n567) & (n1209)));
	assign n1210 = (((!i_32_) & (!i_34_) & (n486) & (!n496)) + ((!i_32_) & (!i_34_) & (n486) & (n496)) + ((!i_32_) & (i_34_) & (n486) & (n496)) + ((i_32_) & (!i_34_) & (!n486) & (!n496)) + ((i_32_) & (!i_34_) & (!n486) & (n496)) + ((i_32_) & (!i_34_) & (n486) & (!n496)) + ((i_32_) & (!i_34_) & (n486) & (n496)) + ((i_32_) & (i_34_) & (!n486) & (n496)) + ((i_32_) & (i_34_) & (n486) & (n496)));
	assign n1214 = (((!i_34_) & (!n649) & (!n974)) + ((!i_34_) & (!n649) & (n974)) + ((!i_34_) & (n649) & (!n974)) + ((!i_34_) & (n649) & (n974)) + ((i_34_) & (!n649) & (n974)) + ((i_34_) & (n649) & (!n974)) + ((i_34_) & (n649) & (n974)));
	assign n1213 = (((!i_30_) & (!n253) & (!n362) & (n1214)) + ((!i_30_) & (!n253) & (n362) & (n1214)) + ((!i_30_) & (n253) & (!n362) & (n1214)) + ((i_30_) & (!n253) & (!n362) & (n1214)) + ((i_30_) & (!n253) & (n362) & (n1214)) + ((i_30_) & (n253) & (!n362) & (n1214)) + ((i_30_) & (n253) & (n362) & (n1214)));
	assign n1215 = (((!n363) & (!n364) & (!n479) & (n498)) + ((!n363) & (!n364) & (n479) & (!n498)) + ((!n363) & (!n364) & (n479) & (n498)) + ((!n363) & (n364) & (!n479) & (n498)) + ((!n363) & (n364) & (n479) & (!n498)) + ((!n363) & (n364) & (n479) & (n498)) + ((n363) & (!n364) & (!n479) & (n498)) + ((n363) & (!n364) & (n479) & (!n498)) + ((n363) & (!n364) & (n479) & (n498)));
	assign n1216 = (((!i_0_) & (n10) & (!n531) & (!n912)) + ((!i_0_) & (n10) & (n531) & (!n912)) + ((i_0_) & (n10) & (!n531) & (!n912)) + ((i_0_) & (n10) & (n531) & (!n912)) + ((i_0_) & (n10) & (n531) & (n912)));
	assign n1222 = (((!n315) & (!n688) & (!n887) & (!n1024)) + ((!n315) & (!n688) & (!n887) & (n1024)) + ((!n315) & (!n688) & (n887) & (!n1024)) + ((!n315) & (!n688) & (n887) & (n1024)) + ((!n315) & (n688) & (!n887) & (!n1024)) + ((!n315) & (n688) & (n887) & (!n1024)) + ((!n315) & (n688) & (n887) & (n1024)) + ((n315) & (!n688) & (!n887) & (!n1024)) + ((n315) & (!n688) & (!n887) & (n1024)) + ((n315) & (!n688) & (n887) & (!n1024)) + ((n315) & (!n688) & (n887) & (n1024)) + ((n315) & (n688) & (!n887) & (!n1024)) + ((n315) & (n688) & (!n887) & (n1024)) + ((n315) & (n688) & (n887) & (!n1024)) + ((n315) & (n688) & (n887) & (n1024)));
	assign n1220 = (((!n668) & (!n995) & (!n1038) & (n1222)) + ((!n668) & (!n995) & (n1038) & (n1222)) + ((!n668) & (n995) & (!n1038) & (n1222)) + ((!n668) & (n995) & (n1038) & (n1222)) + ((n668) & (!n995) & (n1038) & (n1222)) + ((n668) & (n995) & (!n1038) & (n1222)) + ((n668) & (n995) & (n1038) & (n1222)));
	assign n1223 = (((!n494) & (!n874) & (!n1041) & (n1220)) + ((!n494) & (!n874) & (n1041) & (n1220)) + ((!n494) & (n874) & (!n1041) & (n1220)) + ((!n494) & (n874) & (n1041) & (n1220)) + ((n494) & (!n874) & (n1041) & (n1220)) + ((n494) & (n874) & (!n1041) & (n1220)) + ((n494) & (n874) & (n1041) & (n1220)));
	assign n1225 = (((!n315) & (!n572) & (n1038)) + ((!n315) & (n572) & (!n1038)) + ((!n315) & (n572) & (n1038)) + ((n315) & (!n572) & (!n1038)) + ((n315) & (!n572) & (n1038)) + ((n315) & (n572) & (!n1038)) + ((n315) & (n572) & (n1038)));
	assign n1226 = (((!i_14_) & (!n497) & (!n993)) + ((!i_14_) & (!n497) & (n993)) + ((!i_14_) & (n497) & (!n993)) + ((!i_14_) & (n497) & (n993)) + ((i_14_) & (!n497) & (n993)) + ((i_14_) & (n497) & (!n993)) + ((i_14_) & (n497) & (n993)));
	assign n1224 = (((n1225) & (n1226) & (!n873) & (n1041)) + ((n1225) & (n1226) & (n873) & (!n1041)) + ((n1225) & (n1226) & (n873) & (n1041)));
	assign n1228 = (((n455) & (n554)));
	assign n1227 = (((!n864) & (n1042) & (!n1228) & (n813)) + ((!n864) & (n1042) & (n1228) & (!n813)) + ((!n864) & (n1042) & (n1228) & (n813)) + ((n864) & (!n1042) & (!n1228) & (n813)) + ((n864) & (!n1042) & (n1228) & (!n813)) + ((n864) & (!n1042) & (n1228) & (n813)) + ((n864) & (n1042) & (!n1228) & (n813)) + ((n864) & (n1042) & (n1228) & (!n813)) + ((n864) & (n1042) & (n1228) & (n813)));
	assign n1230 = (((!n792) & (!n801) & (!n855)) + ((!n792) & (!n801) & (n855)) + ((!n792) & (n801) & (n855)) + ((n792) & (!n801) & (!n855)) + ((n792) & (!n801) & (n855)) + ((n792) & (n801) & (!n855)) + ((n792) & (n801) & (n855)));
	assign n1229 = (((n1230) & (!n851) & (n170)) + ((n1230) & (n851) & (!n170)) + ((n1230) & (n851) & (n170)));
	assign n1231 = (((!n1276) & (!n170) & (n572)) + ((!n1276) & (n170) & (!n572)) + ((!n1276) & (n170) & (n572)) + ((n1276) & (!n170) & (!n572)) + ((n1276) & (!n170) & (n572)) + ((n1276) & (n170) & (!n572)) + ((n1276) & (n170) & (n572)));
	assign n1232 = (((n681) & (!n809) & (!n810)) + ((n681) & (!n809) & (n810)) + ((n681) & (n809) & (!n810)));
	assign n1237 = (((!n11) & (!n13) & (!n213) & (!n334)) + ((!n11) & (!n13) & (!n213) & (n334)) + ((!n11) & (!n13) & (n213) & (!n334)) + ((!n11) & (!n13) & (n213) & (n334)) + ((!n11) & (n13) & (!n213) & (!n334)) + ((!n11) & (n13) & (!n213) & (n334)) + ((!n11) & (n13) & (n213) & (!n334)) + ((!n11) & (n13) & (n213) & (n334)) + ((n11) & (!n13) & (!n213) & (!n334)) + ((n11) & (!n13) & (!n213) & (n334)) + ((n11) & (!n13) & (n213) & (!n334)) + ((n11) & (!n13) & (n213) & (n334)) + ((n11) & (n13) & (!n213) & (n334)) + ((n11) & (n13) & (n213) & (!n334)) + ((n11) & (n13) & (n213) & (n334)));
	assign n1236 = (((!i_17_) & (!i_21_) & (!n1232) & (n1237)) + ((!i_17_) & (i_21_) & (!n1232) & (n1237)) + ((!i_17_) & (i_21_) & (n1232) & (n1237)) + ((i_17_) & (!i_21_) & (!n1232) & (n1237)) + ((i_17_) & (!i_21_) & (n1232) & (n1237)) + ((i_17_) & (i_21_) & (!n1232) & (n1237)) + ((i_17_) & (i_21_) & (n1232) & (n1237)));
	assign n1238 = (((n1236) & (!i_7_) & (!n973) & (n993)) + ((n1236) & (!i_7_) & (n973) & (!n993)) + ((n1236) & (!i_7_) & (n973) & (n993)) + ((n1236) & (i_7_) & (!n973) & (!n993)) + ((n1236) & (i_7_) & (!n973) & (n993)) + ((n1236) & (i_7_) & (n973) & (!n993)) + ((n1236) & (i_7_) & (n973) & (n993)));
	assign n1239 = (((!i_34_) & (!n253) & (!n823) & (!n827)) + ((!i_34_) & (!n253) & (!n823) & (n827)) + ((!i_34_) & (!n253) & (n823) & (!n827)) + ((!i_34_) & (!n253) & (n823) & (n827)) + ((!i_34_) & (n253) & (!n823) & (n827)) + ((!i_34_) & (n253) & (n823) & (n827)) + ((i_34_) & (!n253) & (n823) & (!n827)) + ((i_34_) & (!n253) & (n823) & (n827)) + ((i_34_) & (n253) & (n823) & (n827)));
	assign n1242 = (((!i_30_) & (!i_36_) & (!n249) & (!n764)) + ((!i_30_) & (!i_36_) & (!n249) & (n764)) + ((!i_30_) & (!i_36_) & (n249) & (!n764)) + ((!i_30_) & (!i_36_) & (n249) & (n764)) + ((!i_30_) & (i_36_) & (!n249) & (n764)) + ((!i_30_) & (i_36_) & (n249) & (!n764)) + ((!i_30_) & (i_36_) & (n249) & (n764)) + ((i_30_) & (!i_36_) & (!n249) & (!n764)) + ((i_30_) & (!i_36_) & (!n249) & (n764)) + ((i_30_) & (!i_36_) & (n249) & (!n764)) + ((i_30_) & (!i_36_) & (n249) & (n764)) + ((i_30_) & (i_36_) & (!n249) & (!n764)) + ((i_30_) & (i_36_) & (!n249) & (n764)) + ((i_30_) & (i_36_) & (n249) & (!n764)) + ((i_30_) & (i_36_) & (n249) & (n764)));
	assign n1241 = (((n953) & (n1011)));
	assign n1244 = (((!i_36_) & (!n13) & (!n192) & (!n364)) + ((!i_36_) & (!n13) & (!n192) & (n364)) + ((!i_36_) & (!n13) & (n192) & (!n364)) + ((!i_36_) & (!n13) & (n192) & (n364)) + ((!i_36_) & (n13) & (!n192) & (!n364)) + ((!i_36_) & (n13) & (!n192) & (n364)) + ((!i_36_) & (n13) & (n192) & (!n364)) + ((!i_36_) & (n13) & (n192) & (n364)) + ((i_36_) & (!n13) & (!n192) & (!n364)) + ((i_36_) & (!n13) & (!n192) & (n364)) + ((i_36_) & (!n13) & (n192) & (!n364)) + ((i_36_) & (!n13) & (n192) & (n364)) + ((i_36_) & (n13) & (!n192) & (!n364)) + ((i_36_) & (n13) & (n192) & (!n364)) + ((i_36_) & (n13) & (n192) & (n364)));
	assign n1243 = (((n614) & (!n793) & (!n951) & (n1244)) + ((n614) & (n793) & (!n951) & (n1244)) + ((n614) & (n793) & (n951) & (n1244)));
	assign n1245 = (((!i_29_) & (n787) & (!n779) & (n812)) + ((!i_29_) & (n787) & (n779) & (!n812)) + ((!i_29_) & (n787) & (n779) & (n812)) + ((i_29_) & (!n787) & (!n779) & (n812)) + ((i_29_) & (!n787) & (n779) & (!n812)) + ((i_29_) & (!n787) & (n779) & (n812)) + ((i_29_) & (n787) & (!n779) & (n812)) + ((i_29_) & (n787) & (n779) & (!n812)) + ((i_29_) & (n787) & (n779) & (n812)));
	assign n1247 = (((!n848) & (!n891) & (!n920)) + ((!n848) & (!n891) & (n920)) + ((!n848) & (n891) & (n920)) + ((n848) & (!n891) & (!n920)) + ((n848) & (!n891) & (n920)) + ((n848) & (n891) & (!n920)) + ((n848) & (n891) & (n920)));
	assign n1246 = (((n1247) & (!n929) & (n558) & (n1019)) + ((n1247) & (n929) & (!n558) & (!n1019)) + ((n1247) & (n929) & (!n558) & (n1019)) + ((n1247) & (n929) & (n558) & (!n1019)) + ((n1247) & (n929) & (n558) & (n1019)));
	assign n1248 = (((n1246) & (!n927) & (n1038)) + ((n1246) & (n927) & (!n1038)) + ((n1246) & (n927) & (n1038)));
	assign n1249 = (((!n362) & (!n872) & (n921) & (!n924)) + ((!n362) & (!n872) & (n921) & (n924)) + ((!n362) & (n872) & (!n921) & (!n924)) + ((!n362) & (n872) & (!n921) & (n924)) + ((!n362) & (n872) & (n921) & (!n924)) + ((!n362) & (n872) & (n921) & (n924)) + ((n362) & (!n872) & (n921) & (n924)) + ((n362) & (n872) & (!n921) & (n924)) + ((n362) & (n872) & (n921) & (n924)));
	assign n1250 = (((!n31) & (!n688) & (n913) & (!n918)) + ((!n31) & (!n688) & (n913) & (n918)) + ((!n31) & (n688) & (n913) & (n918)) + ((n31) & (!n688) & (!n913) & (!n918)) + ((n31) & (!n688) & (!n913) & (n918)) + ((n31) & (!n688) & (n913) & (!n918)) + ((n31) & (!n688) & (n913) & (n918)) + ((n31) & (n688) & (!n913) & (n918)) + ((n31) & (n688) & (n913) & (n918)));
	assign n1251 = (((!i_36_) & (!n852) & (n1039) & (!n1273)) + ((!i_36_) & (!n852) & (n1039) & (n1273)) + ((!i_36_) & (n852) & (!n1039) & (!n1273)) + ((!i_36_) & (n852) & (!n1039) & (n1273)) + ((!i_36_) & (n852) & (n1039) & (!n1273)) + ((!i_36_) & (n852) & (n1039) & (n1273)) + ((i_36_) & (!n852) & (n1039) & (!n1273)) + ((i_36_) & (n852) & (!n1039) & (!n1273)) + ((i_36_) & (n852) & (n1039) & (!n1273)));
	assign n1253 = (((n1251) & (!n664) & (n1245) & (n1243)) + ((n1251) & (n664) & (!n1245) & (!n1243)) + ((n1251) & (n664) & (!n1245) & (n1243)) + ((n1251) & (n664) & (n1245) & (!n1243)) + ((n1251) & (n664) & (n1245) & (n1243)));
	assign n1256 = (((!n608) & (!n501) & (!n654) & (i_29_)) + ((!n608) & (!n501) & (n654) & (!i_29_)) + ((!n608) & (!n501) & (n654) & (i_29_)) + ((!n608) & (n501) & (!n654) & (!i_29_)) + ((!n608) & (n501) & (!n654) & (i_29_)) + ((!n608) & (n501) & (n654) & (!i_29_)) + ((!n608) & (n501) & (n654) & (i_29_)) + ((n608) & (!n501) & (!n654) & (!i_29_)) + ((n608) & (!n501) & (!n654) & (i_29_)) + ((n608) & (!n501) & (n654) & (!i_29_)) + ((n608) & (!n501) & (n654) & (i_29_)) + ((n608) & (n501) & (!n654) & (!i_29_)) + ((n608) & (n501) & (!n654) & (i_29_)) + ((n608) & (n501) & (n654) & (!i_29_)) + ((n608) & (n501) & (n654) & (i_29_)));
	assign n1257 = (((!i_21_) & (!i_36_) & (!n559) & (!n906)) + ((!i_21_) & (!i_36_) & (!n559) & (n906)) + ((!i_21_) & (!i_36_) & (n559) & (!n906)) + ((!i_21_) & (!i_36_) & (n559) & (n906)) + ((!i_21_) & (i_36_) & (!n559) & (n906)) + ((!i_21_) & (i_36_) & (n559) & (!n906)) + ((!i_21_) & (i_36_) & (n559) & (n906)) + ((i_21_) & (!i_36_) & (!n559) & (!n906)) + ((i_21_) & (!i_36_) & (!n559) & (n906)) + ((i_21_) & (!i_36_) & (n559) & (!n906)) + ((i_21_) & (!i_36_) & (n559) & (n906)) + ((i_21_) & (i_36_) & (!n559) & (!n906)) + ((i_21_) & (i_36_) & (!n559) & (n906)) + ((i_21_) & (i_36_) & (n559) & (!n906)) + ((i_21_) & (i_36_) & (n559) & (n906)));
	assign n1258 = (((!i_33_) & (n963)) + ((i_33_) & (!n963)) + ((i_33_) & (n963)));
	assign n1259 = (((!i_13_) & (!n40) & (!n364)) + ((!i_13_) & (n40) & (!n364)) + ((!i_13_) & (n40) & (n364)) + ((i_13_) & (!n40) & (!n364)) + ((i_13_) & (!n40) & (n364)) + ((i_13_) & (n40) & (!n364)) + ((i_13_) & (n40) & (n364)));
	assign n1260 = (((!n558) & (n1018)) + ((n558) & (!n1018)) + ((n558) & (n1018)));
	assign n1261 = (((!n59) & (n763)) + ((n59) & (!n763)) + ((n59) & (n763)));
	assign n1263 = (((!n179) & (!n247) & (!n322)) + ((!n179) & (n247) & (!n322)) + ((!n179) & (n247) & (n322)) + ((n179) & (!n247) & (!n322)) + ((n179) & (!n247) & (n322)) + ((n179) & (n247) & (!n322)) + ((n179) & (n247) & (n322)));
	assign n1264 = (((!i_24_) & (!i_28_) & (n289)) + ((!i_24_) & (i_28_) & (!n289)) + ((!i_24_) & (i_28_) & (n289)) + ((i_24_) & (!i_28_) & (!n289)) + ((i_24_) & (!i_28_) & (n289)) + ((i_24_) & (i_28_) & (!n289)) + ((i_24_) & (i_28_) & (n289)));
	assign n1268 = (((!i_0_) & (!n500) & (!n511) & (!n800)) + ((!i_0_) & (!n500) & (n511) & (!n800)) + ((!i_0_) & (!n500) & (n511) & (n800)) + ((!i_0_) & (n500) & (!n511) & (!n800)) + ((!i_0_) & (n500) & (!n511) & (n800)) + ((!i_0_) & (n500) & (n511) & (!n800)) + ((!i_0_) & (n500) & (n511) & (n800)) + ((i_0_) & (!n500) & (!n511) & (!n800)) + ((i_0_) & (!n500) & (!n511) & (n800)) + ((i_0_) & (!n500) & (n511) & (!n800)) + ((i_0_) & (!n500) & (n511) & (n800)) + ((i_0_) & (n500) & (!n511) & (!n800)) + ((i_0_) & (n500) & (!n511) & (n800)) + ((i_0_) & (n500) & (n511) & (!n800)) + ((i_0_) & (n500) & (n511) & (n800)));
	assign n1272 = (((n482) & (n1029)));
	assign n1273 = (((!n834) & (!n837) & (!n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (!n843) & (n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (!n840) & (n843) & (n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (!n843) & (n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (!n837) & (n840) & (n843) & (n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (!n843) & (n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (!n840) & (n843) & (n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (!n843) & (n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((!n834) & (n837) & (n840) & (n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((!n834) & (n837) & (n840) & (n843) & (n845) & (n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (!n843) & (n845) & (n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (!n840) & (n843) & (n845) & (n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (!n843) & (n845) & (n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (!n837) & (n840) & (n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (!n837) & (n840) & (n843) & (n845) & (n847) & (n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (!n843) & (n845) & (n847) & (n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (!n840) & (n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (!n840) & (n843) & (n845) & (n847) & (n1238) & (n1239)) + ((n834) & (n837) & (n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (!n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (n840) & (!n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (!n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (n837) & (n840) & (!n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (!n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (n840) & (!n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (!n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((n834) & (n837) & (n840) & (!n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (!n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (n840) & (!n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (!n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (n837) & (n840) & (!n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (!n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (n840) & (!n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (!n843) & (n845) & (n847) & (n1238) & (n1239)) + ((n834) & (n837) & (n840) & (n843) & (!n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (n843) & (!n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (n840) & (n843) & (!n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (n843) & (!n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (n837) & (n840) & (n843) & (!n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (n843) & (!n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (n840) & (n843) & (!n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (n843) & (!n845) & (n847) & (n1238) & (n1239)) + ((n834) & (n837) & (n840) & (n843) & (n845) & (!n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (n843) & (n845) & (!n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (n840) & (n843) & (n845) & (!n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (n843) & (n845) & (!n847) & (n1238) & (n1239)) + ((n834) & (n837) & (n840) & (n843) & (n845) & (n847) & (!n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (n843) & (n845) & (n847) & (!n1238) & (n1239)) + ((n834) & (n837) & (n840) & (n843) & (n845) & (n847) & (n1238) & (!n1239)) + ((n834) & (n837) & (n840) & (n843) & (n845) & (n847) & (n1238) & (n1239)));
	assign n1276 = (((n646) & (n1022)));
	assign n1279 = (((!n163) & (n290) & (n670)));
	assign n1280 = (((!i_23_) & (!n10) & (!n522) & (!n901)) + ((!i_23_) & (!n10) & (!n522) & (n901)) + ((!i_23_) & (!n10) & (n522) & (!n901)) + ((!i_23_) & (!n10) & (n522) & (n901)) + ((!i_23_) & (n10) & (!n522) & (n901)) + ((!i_23_) & (n10) & (n522) & (!n901)) + ((!i_23_) & (n10) & (n522) & (n901)) + ((i_23_) & (!n10) & (!n522) & (!n901)) + ((i_23_) & (!n10) & (!n522) & (n901)) + ((i_23_) & (!n10) & (n522) & (!n901)) + ((i_23_) & (!n10) & (n522) & (n901)) + ((i_23_) & (n10) & (!n522) & (!n901)) + ((i_23_) & (n10) & (!n522) & (n901)) + ((i_23_) & (n10) & (n522) & (!n901)) + ((i_23_) & (n10) & (n522) & (n901)));
	assign n1281 = (((i_0_) & (!i_12_) & (n10) & (n531) & (n801)));

endmodule