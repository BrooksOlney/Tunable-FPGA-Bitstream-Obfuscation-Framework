module apex4x5xv (i_7_, i_8_, i_5_, i_6_, i_3_, i_4_, i_1_, i_2_, i_0_, o_1_, o_2_, o_12_, o_11_, o_14_, o_13_, o_16_, o_15_, o_18_, o_17_, o_10_, o_9_, o_7_, o_8_, o_5_, o_6_, o_3_, o_4_);

	input i_7_;
	input i_8_;
	input i_5_;
	input i_6_;
	input i_3_;
	input i_4_;
	input i_1_;
	input i_2_;
	input i_0_;
	output o_1_;
	output o_2_;
	output o_12_;
	output o_11_;
	output o_14_;
	output o_13_;
	output o_16_;
	output o_15_;
	output o_18_;
	output o_17_;
	output o_10_;
	output o_9_;
	output o_7_;
	output o_8_;
	output o_5_;
	output o_6_;
	output o_3_;
	output o_4_;

	wire [963 : 0] sk /* synthesis noprune */;

	lut_sub lut_3 ({sk[0], x4869x, x4838x, x4839x, x4865x}, o_1_);
	defparam lut_3.LUT_SIZE = 5;
	defparam lut_3.mask = 32'h33ff7fff;

	lut_sub lut_8 ({sk[1], x4991x, x4992x}, o_2_);
	defparam lut_8.LUT_SIZE = 3;
	defparam lut_8.mask = 8'h37;

	lut_sub lut_11 ({sk[2], x5048x, x5010x, x5011x, x5029x, x5030x}, o_12_);
	defparam lut_11.LUT_SIZE = 6;
	defparam lut_11.mask = 64'h05ffffff7fffffff;

	lut_sub lut_17 ({sk[3], n_n722, n_n724, x5108x, x6347x}, o_11_);
	defparam lut_17.LUT_SIZE = 5;
	defparam lut_17.mask = 32'h33ffbfff;

	lut_sub lut_22 ({sk[4], x5168x, x5139x, x5140x, x5164x, x5165x}, o_14_);
	defparam lut_22.LUT_SIZE = 6;
	defparam lut_22.mask = 64'h05ffffff7fffffff;

	lut_sub lut_28 ({sk[5], x5221x, x5218x, x5219x}, o_13_);
	defparam lut_28.LUT_SIZE = 4;
	defparam lut_28.mask = 16'h0f7f;

	lut_sub lut_32 ({sk[6], x5232x, x178x, x258x, x310x, x5230x}, o_16_);
	defparam lut_32.LUT_SIZE = 6;
	defparam lut_32.mask = 64'h05ffffff7fffffff;

	lut_sub lut_38 ({sk[7], x5250x, x310x, x188x, x114x, x5246x}, o_15_);
	defparam lut_38.LUT_SIZE = 6;
	defparam lut_38.mask = 64'h05ffffff7fffffff;

	lut_sub lut_44 ({sk[8], x5265x, x5260x, x5261x}, o_18_);
	defparam lut_44.LUT_SIZE = 4;
	defparam lut_44.mask = 16'h0f7f;

	lut_sub lut_48 ({sk[9], x5270x, x187x, x259x, x294x, x261x}, o_17_);
	defparam lut_48.LUT_SIZE = 6;
	defparam lut_48.mask = 64'h05ffffff7fffffff;

	lut_sub lut_54 ({sk[10], x5373x, x5315x, x5316x, x5369x, x5370x}, o_10_);
	defparam lut_54.LUT_SIZE = 6;
	defparam lut_54.mask = 64'h05ffffff7fffffff;

	lut_sub lut_60 ({sk[11], x5490x, x5485x, x5486x, x5488x}, o_9_);
	defparam lut_60.LUT_SIZE = 5;
	defparam lut_60.mask = 32'h33ff7fff;

	lut_sub lut_65 ({sk[12], n_n444, n_n450, x5586x, x5587x, x5588x}, o_7_);
	defparam lut_65.LUT_SIZE = 6;
	defparam lut_65.mask = 64'h05ffffff7fffffff;

	lut_sub lut_71 ({sk[13], x5685x, n_n517, x5654x, x5655x, x5656x}, o_8_);
	defparam lut_71.LUT_SIZE = 6;
	defparam lut_71.mask = 64'h05ffffff7fffffff;

	lut_sub lut_77 ({sk[14], x5781x, x5732x, n_n305, x5731x}, o_5_);
	defparam lut_77.LUT_SIZE = 5;
	defparam lut_77.mask = 32'h33ff7fff;

	lut_sub lut_82 ({sk[15], x5877x, n_n377, x5818x, x5819x, x5820x}, o_6_);
	defparam lut_82.LUT_SIZE = 6;
	defparam lut_82.mask = 64'h05ffffff7fffffff;

	lut_sub lut_88 ({sk[16], x5942x, x5937x, x5938x}, o_3_);
	defparam lut_88.LUT_SIZE = 4;
	defparam lut_88.mask = 16'h0f7f;

	lut_sub lut_92 ({sk[17], x6028x, x6029x}, o_4_);
	defparam lut_92.LUT_SIZE = 3;
	defparam lut_92.mask = 8'h37;

	lut_sub lut_95 ({sk[18], x4855x, x4856x, x4861x, x4862x, x4864x}, x4869x);
	defparam lut_95.LUT_SIZE = 6;
	defparam lut_95.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_101 ({sk[19], n_n78, x42x, n_n1120, x355x, n_n1156}, x4838x);
	defparam lut_101.LUT_SIZE = 6;
	defparam lut_101.mask = 64'h7fff7fff7f7f7fff;

	lut_sub lut_106 ({sk[20], i_6_, n_n86, x42x, n_n1021, x4837x}, x4839x);
	defparam lut_106.LUT_SIZE = 6;
	defparam lut_106.mask = 64'h7fff7fff7777777f;

	lut_sub lut_110 ({sk[21], n_n80, x337x, x1589x, x4848x, x4860x}, x4865x);
	defparam lut_110.LUT_SIZE = 6;
	defparam lut_110.mask = 64'h7fff7fff7f7f7fff;

	lut_sub lut_115 ({sk[22], x4928x, x4929x, x232x, x4984x, x4987x}, x4991x);
	defparam lut_115.LUT_SIZE = 6;
	defparam lut_115.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_121 ({sk[23], n_n131, x4919x, x4920x, x4985x, x4986x}, x4992x);
	defparam lut_121.LUT_SIZE = 6;
	defparam lut_121.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_127 ({sk[24], x5038x, x5039x, x5040x, x5041x, x5046x}, x5048x);
	defparam lut_127.LUT_SIZE = 6;
	defparam lut_127.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_133 ({sk[25], n_n73, x21x, x256x, x299x, x5006x}, x5010x);
	defparam lut_133.LUT_SIZE = 6;
	defparam lut_133.mask = 64'h7fff7fff7f7f7fff;

	lut_sub lut_138 ({sk[26], x190x, x265x, x5003x, x5004x, x5005x}, x5011x);
	defparam lut_138.LUT_SIZE = 6;
	defparam lut_138.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_144 ({sk[27], x135x, n_n949, x97x, x204x, x5025x}, x5029x);
	defparam lut_144.LUT_SIZE = 6;
	defparam lut_144.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_150 ({sk[28], x195x, x151x, x5021x, x5023x, x5024x}, x5030x);
	defparam lut_150.LUT_SIZE = 6;
	defparam lut_150.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_156 ({sk[29], x5060x, x5061x, x5062x, x5063x, x5064x}, n_n722);
	defparam lut_156.LUT_SIZE = 6;
	defparam lut_156.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_162 ({sk[30], x5076x, x5077x, x5078x, x5079x}, n_n724);
	defparam lut_162.LUT_SIZE = 5;
	defparam lut_162.mask = 32'h33ff7fff;

	lut_sub lut_167 ({sk[31], n_n1324, n_n1092, x5087x, x5099x, x5104x}, x5108x);
	defparam lut_167.LUT_SIZE = 6;
	defparam lut_167.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_173 ({sk[32], x257x, x5093x, x5100x, x5101x, x5103x}, x6347x);
	defparam lut_173.LUT_SIZE = 6;
	defparam lut_173.mask = 64'h7fff7fff80000000;

	lut_sub lut_175 ({sk[33], n_n846, x5154x, x5155x, x5156x, x5157x}, x5168x);
	defparam lut_175.LUT_SIZE = 6;
	defparam lut_175.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_181 ({sk[34], n_n38, x52x, x306x, x1480x, x5135x}, x5139x);
	defparam lut_181.LUT_SIZE = 6;
	defparam lut_181.mask = 64'h7fff7fff7f7f7fff;

	lut_sub lut_186 ({sk[35], x141x, x279x, x5131x, x5133x, x5134x}, x5140x);
	defparam lut_186.LUT_SIZE = 6;
	defparam lut_186.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_192 ({sk[36], x64x, n_n82, x342x, x5148x, x5159x}, x5164x);
	defparam lut_192.LUT_SIZE = 6;
	defparam lut_192.mask = 64'h7fff7fff7f7f7fff;

	lut_sub lut_197 ({sk[37], x123x, x183x, x5150x, x5151x, x5152x}, x5165x);
	defparam lut_197.LUT_SIZE = 6;
	defparam lut_197.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_203 ({sk[38], x5185x, x5186x, x5202x, x5203x}, x5221x);
	defparam lut_203.LUT_SIZE = 5;
	defparam lut_203.mask = 32'h33ff7fff;

	lut_sub lut_208 ({sk[39], x178x, x1413x, x1414x, x5208x, x5214x}, x5218x);
	defparam lut_208.LUT_SIZE = 6;
	defparam lut_208.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_214 ({sk[40], x1285x, x186x, x5217x, x6355x}, x5219x);
	defparam lut_214.LUT_SIZE = 5;
	defparam lut_214.mask = 32'h33ffbfff;

	lut_sub lut_219 ({sk[41], n_n1369, n_n1176, x187x, x259x, x294x}, x5232x);
	defparam lut_219.LUT_SIZE = 6;
	defparam lut_219.mask = 64'h7fff7fff7fffffff;

	lut_sub lut_225 ({sk[42], i_7_, i_8_, i_6_, x76x, x43x}, x178x);
	defparam lut_225.LUT_SIZE = 6;
	defparam lut_225.mask = 64'h7fff7fff50030000;

	lut_sub lut_228 ({sk[43], n_n78, n_n91, n_n92, n_n74, n_n90}, x258x);
	defparam lut_228.LUT_SIZE = 6;
	defparam lut_228.mask = 64'h7fff7fff00110515;

	lut_sub lut_231 ({sk[44], n_n1297, n_n1283, n_n1312, x326x}, x310x);
	defparam lut_231.LUT_SIZE = 5;
	defparam lut_231.mask = 32'h33ff7fff;

	lut_sub lut_236 ({sk[45], n_n38, n_n93, x43x, n_n1074, n_n1294}, x5230x);
	defparam lut_236.LUT_SIZE = 6;
	defparam lut_236.mask = 64'h7fff7fff777f7f7f;

	lut_sub lut_241 ({sk[46], x136x, x230x, x5242x, x5248x}, x5250x);
	defparam lut_241.LUT_SIZE = 5;
	defparam lut_241.mask = 32'h33ff7fff;

	lut_sub lut_246 ({sk[47], i_3_, n_n101, x325x, n_n90, n_n1047}, x188x);
	defparam lut_246.LUT_SIZE = 6;
	defparam lut_246.mask = 64'h0055ffff55555557;

	lut_sub lut_249 ({sk[48], i_3_, n_n78, n_n94, x325x, n_n1042}, x114x);
	defparam lut_249.LUT_SIZE = 6;
	defparam lut_249.mask = 64'h0055ffff55555557;

	lut_sub lut_252 ({sk[49], n_n1281, n_n1279, x258x, x259x, x294x}, x5246x);
	defparam lut_252.LUT_SIZE = 6;
	defparam lut_252.mask = 64'h0055ffff7fffffff;

	lut_sub lut_258 ({sk[50], x230x, x261x, x5259x, x5262x}, x5265x);
	defparam lut_258.LUT_SIZE = 5;
	defparam lut_258.mask = 32'h0f7f7fff;

	lut_sub lut_263 ({sk[51], n_n1294, n_n1169, n_n942, n_n1057}, x5260x);
	defparam lut_263.LUT_SIZE = 5;
	defparam lut_263.mask = 32'h0f7f7fff;

	lut_sub lut_268 ({sk[52], n_n101, x43x, n_n1125, n_n1128, n_n1286}, x5261x);
	defparam lut_268.LUT_SIZE = 6;
	defparam lut_268.mask = 64'h0055ffff7f7f7fff;

	lut_sub lut_273 ({sk[53], n_n63, x49x, n_n1176, x248x, n_n1283}, x5270x);
	defparam lut_273.LUT_SIZE = 6;
	defparam lut_273.mask = 64'h0055ffff7f7f7fff;

	lut_sub lut_278 ({sk[54], i_3_, x341x, n_n95, x36x, x31x}, x187x);
	defparam lut_278.LUT_SIZE = 6;
	defparam lut_278.mask = 64'h0055ffff03030357;

	lut_sub lut_281 ({sk[55], i_5_, n_n101, x54x, n_n90, n_n1132}, x259x);
	defparam lut_281.LUT_SIZE = 6;
	defparam lut_281.mask = 64'h0055ffff55575555;

	lut_sub lut_284 ({sk[56], i_1_, i_2_, i_0_, x131x, x5012x}, x294x);
	defparam lut_284.LUT_SIZE = 6;
	defparam lut_284.mask = 64'h00ff33fff0700000;

	lut_sub lut_288 ({sk[57], i_7_, i_8_, i_6_, x39x, n_n941}, x261x);
	defparam lut_288.LUT_SIZE = 6;
	defparam lut_288.mask = 64'h00ff33ff55555575;

	lut_sub lut_291 ({sk[58], x5331x, x5332x, x5333x, x5334x, x5371x}, x5373x);
	defparam lut_291.LUT_SIZE = 6;
	defparam lut_291.mask = 64'h00ff33ff7fffffff;

	lut_sub lut_297 ({sk[59], x5273x, x5274x, x5306x, x5307x}, x5315x);
	defparam lut_297.LUT_SIZE = 5;
	defparam lut_297.mask = 32'h3f3f7fff;

	lut_sub lut_302 ({sk[60], x5298x, x5309x, x5310x, x6345x}, x5316x);
	defparam lut_302.LUT_SIZE = 5;
	defparam lut_302.mask = 32'h3f3fbfff;

	lut_sub lut_307 ({sk[61], n_n1082, x1487x, x90x, x298x, x5364x}, x5369x);
	defparam lut_307.LUT_SIZE = 6;
	defparam lut_307.mask = 64'h00ff33ff7fffffff;

	lut_sub lut_313 ({sk[62], n_n958, x5358x, x5359x, x6344x, x6351x}, x5370x);
	defparam lut_313.LUT_SIZE = 6;
	defparam lut_313.mask = 64'h00ff33ffefffffff;

	lut_sub lut_319 ({sk[63], x5388x, x5389x, x5403x, x5404x, x5484x}, x5490x);
	defparam lut_319.LUT_SIZE = 6;
	defparam lut_319.mask = 64'h00ffffff7fffffff;

	lut_sub lut_325 ({sk[64], x5450x, x335x, x1440x, x5446x, x5482x}, x5485x);
	defparam lut_325.LUT_SIZE = 6;
	defparam lut_325.mask = 64'h00ffffff7fffffff;

	lut_sub lut_331 ({sk[65], x5454x, x263x, x91x, x5478x, x5479x}, x5486x);
	defparam lut_331.LUT_SIZE = 6;
	defparam lut_331.mask = 64'h00ffffff7fffffff;

	lut_sub lut_337 ({sk[66], x5421x, x5422x, x5440x, x5441x}, x5488x);
	defparam lut_337.LUT_SIZE = 5;
	defparam lut_337.mask = 32'h0f0f7fff;

	lut_sub lut_342 ({sk[67], x5539x, x5513x, x5508x, x5509x, x5538x}, n_n444);
	defparam lut_342.LUT_SIZE = 6;
	defparam lut_342.mask = 64'h00ffffff7fffffff;

	lut_sub lut_348 ({sk[68], x5550x, x5551x, x5552x, x5553x, x5554x}, n_n450);
	defparam lut_348.LUT_SIZE = 6;
	defparam lut_348.mask = 64'h00ffffff7fffffff;

	lut_sub lut_354 ({sk[69], x204x, x263x, x5571x, x5580x}, x5586x);
	defparam lut_354.LUT_SIZE = 5;
	defparam lut_354.mask = 32'h0f0f7fff;

	lut_sub lut_359 ({sk[70], x5573x, x5574x, x5575x, x5576x}, x5587x);
	defparam lut_359.LUT_SIZE = 5;
	defparam lut_359.mask = 32'h0f0f7fff;

	lut_sub lut_364 ({sk[71], x168x, x5568x, x5579x, x6358x}, x5588x);
	defparam lut_364.LUT_SIZE = 5;
	defparam lut_364.mask = 32'h0f0fbfff;

	lut_sub lut_369 ({sk[72], n_n514, x5676x, x5677x, x5680x, x5682x}, x5685x);
	defparam lut_369.LUT_SIZE = 6;
	defparam lut_369.mask = 64'h00ffffff7fffffff;

	lut_sub lut_375 ({sk[73], x5616x, x5617x, x5618x, x5619x, x5620x}, n_n517);
	defparam lut_375.LUT_SIZE = 6;
	defparam lut_375.mask = 64'h00ffffff7fffffff;

	lut_sub lut_381 ({sk[74], x94x, x195x, x223x, x101x, x5648x}, x5654x);
	defparam lut_381.LUT_SIZE = 6;
	defparam lut_381.mask = 64'h00ffffff7fffffff;

	lut_sub lut_387 ({sk[75], x5641x, x5642x, x5643x, x5644x}, x5655x);
	defparam lut_387.LUT_SIZE = 5;
	defparam lut_387.mask = 32'h0f0f7fff;

	lut_sub lut_392 ({sk[76], x97x, x125x, x5645x, x5646x, x6340x}, x5656x);
	defparam lut_392.LUT_SIZE = 6;
	defparam lut_392.mask = 64'h00ffffffbfffffff;

	lut_sub lut_398 ({sk[77], n_n308, x5773x, x5774x, x5776x, x5778x}, x5781x);
	defparam lut_398.LUT_SIZE = 6;
	defparam lut_398.mask = 64'h00ffffff7fffffff;

	lut_sub lut_404 ({sk[78], n_n1160, x617x, x5717x, x5726x, x5729x}, x5732x);
	defparam lut_404.LUT_SIZE = 6;
	defparam lut_404.mask = 64'h00ffffff7fffffff;

	lut_sub lut_410 ({sk[79], x5699x, x5700x, x5703x, x5704x, x5706x}, n_n305);
	defparam lut_410.LUT_SIZE = 6;
	defparam lut_410.mask = 64'h00ffffff7fffffff;

	lut_sub lut_416 ({sk[80], x160x, x166x, x281x, x121x, x5727x}, x5731x);
	defparam lut_416.LUT_SIZE = 6;
	defparam lut_416.mask = 64'h00ffffff7fffffff;

	lut_sub lut_422 ({sk[81], n_n376, x5869x, x5870x, x5872x, x5874x}, x5877x);
	defparam lut_422.LUT_SIZE = 6;
	defparam lut_422.mask = 64'h00ffffff7fffffff;

	lut_sub lut_428 ({sk[82], x5791x, x5792x, x5793x, x6333x}, n_n377);
	defparam lut_428.LUT_SIZE = 5;
	defparam lut_428.mask = 32'h0f0fbfff;

	lut_sub lut_433 ({sk[83], x215x, x153x, x103x, n_n959, x5814x}, x5818x);
	defparam lut_433.LUT_SIZE = 6;
	defparam lut_433.mask = 64'h00ffffff7fffffff;

	lut_sub lut_439 ({sk[84], n_n944, n_n939, x5399x, x5808x, x6357x}, x5819x);
	defparam lut_439.LUT_SIZE = 6;
	defparam lut_439.mask = 64'h00ffffffbfffffff;

	lut_sub lut_445 ({sk[85], x303x, n_n652, x5809x, x5810x, x5812x}, x5820x);
	defparam lut_445.LUT_SIZE = 6;
	defparam lut_445.mask = 64'h00ffffff7fffffff;

	lut_sub lut_451 ({sk[86], x5896x, x5897x, x5934x, x5935x, x5936x}, x5942x);
	defparam lut_451.LUT_SIZE = 6;
	defparam lut_451.mask = 64'h00ffffff7fffffff;

	lut_sub lut_457 ({sk[87], x103x, x5901x, n_n984, x5899x, x5933x}, x5937x);
	defparam lut_457.LUT_SIZE = 6;
	defparam lut_457.mask = 64'h00ffffff7fffffff;

	lut_sub lut_463 ({sk[88], x153x, x5904x, x5907x, x5908x, n_n952}, x5938x);
	defparam lut_463.LUT_SIZE = 6;
	defparam lut_463.mask = 64'h00ffffff7fffffff;

	lut_sub lut_469 ({sk[89], x5953x, x5954x, x5955x, x5956x, x6026x}, x6028x);
	defparam lut_469.LUT_SIZE = 6;
	defparam lut_469.mask = 64'h00ffffff7fffffff;

	lut_sub lut_475 ({sk[90], x5987x, x5985x, x5986x, x6024x, x6025x}, x6029x);
	defparam lut_475.LUT_SIZE = 6;
	defparam lut_475.mask = 64'h00ffffff7fffffff;

	lut_sub lut_481 ({sk[91], x57x, n_n92, x113x, n_n95, x132x}, x4855x);
	defparam lut_481.LUT_SIZE = 6;
	defparam lut_481.mask = 64'h00ffffff0f5f3f7f;

	lut_sub lut_485 ({sk[92], x27x, n_n63, x208x, n_n95, x34x}, x4856x);
	defparam lut_485.LUT_SIZE = 6;
	defparam lut_485.mask = 64'h00ffffff0f5f3f7f;

	lut_sub lut_489 ({sk[93], n_n101, n_n91, n_n83, n_n102, x4852x}, x4861x);
	defparam lut_489.LUT_SIZE = 6;
	defparam lut_489.mask = 64'h00ffffff55575757;

	lut_sub lut_493 ({sk[94], n_n58, x26x, x39x, x87x, x104x}, x4862x);
	defparam lut_493.LUT_SIZE = 6;
	defparam lut_493.mask = 64'h00ffffff77777fff;

	lut_sub lut_498 ({sk[95], n_n91, x76x, n_n1185, x227x, x4858x}, x4864x);
	defparam lut_498.LUT_SIZE = 6;
	defparam lut_498.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_503 ({sk[96], n_n91, x49x, x111x, x41x, x136x}, x4928x);
	defparam lut_503.LUT_SIZE = 6;
	defparam lut_503.mask = 64'h00ffffff575757ff;

	lut_sub lut_507 ({sk[97], x27x, x26x, n_n63, n_n82, x4927x}, x4929x);
	defparam lut_507.LUT_SIZE = 6;
	defparam lut_507.mask = 64'h00ffffff55775f7f;

	lut_sub lut_511 ({sk[98], i_4_, n_n93, n_n67, x1479x, x1480x}, x232x);
	defparam lut_511.LUT_SIZE = 6;
	defparam lut_511.mask = 64'h00ffffff777f7777;

	lut_sub lut_515 ({sk[99], x4971x, x4972x, x4973x, x4974x}, x4984x);
	defparam lut_515.LUT_SIZE = 5;
	defparam lut_515.mask = 32'h0f0f7fff;

	lut_sub lut_520 ({sk[100], x4943x, x4950x, x4951x, n_n1215, x121x}, x4987x);
	defparam lut_520.LUT_SIZE = 6;
	defparam lut_520.mask = 64'h00ffffff7fffffff;

	lut_sub lut_526 ({sk[101], x4899x, x4891x, x4892x, x4898x}, n_n131);
	defparam lut_526.LUT_SIZE = 5;
	defparam lut_526.mask = 32'h0f0f7fff;

	lut_sub lut_531 ({sk[102], x298x, x292x, n_n882, x4910x}, x4919x);
	defparam lut_531.LUT_SIZE = 5;
	defparam lut_531.mask = 32'h0f0f7fff;

	lut_sub lut_536 ({sk[103], x4913x, x4914x, x4917x}, x4920x);
	defparam lut_536.LUT_SIZE = 4;
	defparam lut_536.mask = 16'h777f;

	lut_sub lut_540 ({sk[104], x4975x, x4976x, x4982x}, x4985x);
	defparam lut_540.LUT_SIZE = 4;
	defparam lut_540.mask = 16'h777f;

	lut_sub lut_544 ({sk[105], n_n137, x4936x, x231x, x4935x}, x4986x);
	defparam lut_544.LUT_SIZE = 5;
	defparam lut_544.mask = 32'h0f0f7fff;

	lut_sub lut_549 ({sk[106], x32x, n_n77, x346x, x1413x, x1414x}, x5038x);
	defparam lut_549.LUT_SIZE = 6;
	defparam lut_549.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_554 ({sk[107], i_5_, x54x, x343x, x255x, x48x}, x5039x);
	defparam lut_554.LUT_SIZE = 6;
	defparam lut_554.mask = 64'h00ffffff3f3f3f7f;

	lut_sub lut_558 ({sk[108], n_n78, n_n63, x49x, n_n1204, n_n1369}, x5040x);
	defparam lut_558.LUT_SIZE = 6;
	defparam lut_558.mask = 64'h00ffffff777f7f7f;

	lut_sub lut_563 ({sk[109], n_n58, n_n78, x25x, x53x, x5035x}, x5041x);
	defparam lut_563.LUT_SIZE = 6;
	defparam lut_563.mask = 64'h00ffffff55775f7f;

	lut_sub lut_567 ({sk[110], x87x, x61x, x231x, x301x, x5037x}, x5046x);
	defparam lut_567.LUT_SIZE = 6;
	defparam lut_567.mask = 64'h00ffffff7fffffff;

	lut_sub lut_573 ({sk[111], n_n882, x296x, x5121x, x5123x, x5124x}, n_n846);
	defparam lut_573.LUT_SIZE = 6;
	defparam lut_573.mask = 64'h00ffffff7fffffff;

	lut_sub lut_579 ({sk[112], i_5_, x54x, x1285x, x186x, x31x}, x5154x);
	defparam lut_579.LUT_SIZE = 6;
	defparam lut_579.mask = 64'h00ffffff3f3f3f7f;

	lut_sub lut_583 ({sk[113], i_7_, i_6_, x34x, x206x, n_n1215}, x5155x);
	defparam lut_583.LUT_SIZE = 6;
	defparam lut_583.mask = 64'h00ffffff7777777f;

	lut_sub lut_587 ({sk[114], i_1_, n_n86, n_n1324, n_n1369, x72x}, x5156x);
	defparam lut_587.LUT_SIZE = 6;
	defparam lut_587.mask = 64'h00ffffff3f7f3f3f;

	lut_sub lut_591 ({sk[115], n_n63, x49x, n_n1193, n_n1330, n_n1267}, x5157x);
	defparam lut_591.LUT_SIZE = 6;
	defparam lut_591.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_596 ({sk[116], x306x, x5176x, x5181x}, x5185x);
	defparam lut_596.LUT_SIZE = 4;
	defparam lut_596.mask = 16'h777f;

	lut_sub lut_600 ({sk[117], x254x, x88x, x5178x, x5179x, x5180x}, x5186x);
	defparam lut_600.LUT_SIZE = 6;
	defparam lut_600.mask = 64'h00ffffff7fffffff;

	lut_sub lut_606 ({sk[118], x125x, x5193x, x5198x}, x5202x);
	defparam lut_606.LUT_SIZE = 4;
	defparam lut_606.mask = 16'h777f;

	lut_sub lut_610 ({sk[119], x5196x, x5197x, x5200x}, x5203x);
	defparam lut_610.LUT_SIZE = 4;
	defparam lut_610.mask = 16'h777f;

	lut_sub lut_614 ({sk[120], i_7_, i_8_, i_5_, i_6_, x351x}, n_n1369);
	defparam lut_614.LUT_SIZE = 6;
	defparam lut_614.mask = 64'h00ffffff00400000;

	lut_sub lut_616 ({sk[121], i_1_, i_2_, i_0_, n_n91, n_n74}, n_n1176);
	defparam lut_616.LUT_SIZE = 6;
	defparam lut_616.mask = 64'h00ffffff00001000;

	lut_sub lut_618 ({sk[122], i_5_, i_3_, i_4_, x37x, n_n1330}, x136x);
	defparam lut_618.LUT_SIZE = 6;
	defparam lut_618.mask = 64'h00ffffff55555575;

	lut_sub lut_621 ({sk[123], i_7_, i_8_, i_6_, x49x, x333x}, x230x);
	defparam lut_621.LUT_SIZE = 6;
	defparam lut_621.mask = 64'h00ffffff55557555;

	lut_sub lut_624 ({sk[124], n_n93, n_n102, n_n1369, n_n90, x278x}, x5242x);
	defparam lut_624.LUT_SIZE = 6;
	defparam lut_624.mask = 64'h00ffffff5f5f5f7f;

	lut_sub lut_628 ({sk[125], n_n1259, n_n1032, n_n1169, n_n942, x5244x}, x5248x);
	defparam lut_628.LUT_SIZE = 6;
	defparam lut_628.mask = 64'h00ffffff7fffffff;

	lut_sub lut_634 ({sk[126], i_1_, n_n86, n_n1324, x72x, n_n1074}, x5259x);
	defparam lut_634.LUT_SIZE = 6;
	defparam lut_634.mask = 64'h00ffffff5f7f5f5f;

	lut_sub lut_638 ({sk[127], x136x, x114x, x189x, n_n1046, n_n1047}, x5262x);
	defparam lut_638.LUT_SIZE = 6;
	defparam lut_638.mask = 64'h00ffffff7fffffff;

	lut_sub lut_644 ({sk[128], i_7_, i_8_, i_6_}, n_n63);
	defparam lut_644.LUT_SIZE = 4;
	defparam lut_644.mask = 16'h7720;

	lut_sub lut_646 ({sk[129], i_5_, i_3_, i_4_, i_0_, x75x}, x49x);
	defparam lut_646.LUT_SIZE = 6;
	defparam lut_646.mask = 64'h00ffffff00000040;

	lut_sub lut_648 ({sk[130], i_1_, i_2_, i_0_, n_n95, n_n77}, x248x);
	defparam lut_648.LUT_SIZE = 6;
	defparam lut_648.mask = 64'h00ffffff00001000;

	lut_sub lut_650 ({sk[131], i_5_, i_3_, i_4_, n_n91, n_n90}, n_n1283);
	defparam lut_650.LUT_SIZE = 6;
	defparam lut_650.mask = 64'h00ffffff00001000;

	lut_sub lut_652 ({sk[132], x57x, n_n63, n_n1047, n_n1028, n_n1018}, x5331x);
	defparam lut_652.LUT_SIZE = 6;
	defparam lut_652.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_657 ({sk[133], n_n1032, n_n1040, n_n1011, x59x, x1085x}, x5332x);
	defparam lut_657.LUT_SIZE = 6;
	defparam lut_657.mask = 64'h00ffffff7fffffff;

	lut_sub lut_663 ({sk[134], x201x, x164x, x288x, x203x}, x5333x);
	defparam lut_663.LUT_SIZE = 5;
	defparam lut_663.mask = 32'h0f0f7fff;

	lut_sub lut_668 ({sk[135], n_n999, n_n1009, x156x, x5321x, x5322x}, x5334x);
	defparam lut_668.LUT_SIZE = 6;
	defparam lut_668.mask = 64'h00ffffff7fffffff;

	lut_sub lut_674 ({sk[136], x232x, x257x, x168x, x5360x, x5362x}, x5371x);
	defparam lut_674.LUT_SIZE = 6;
	defparam lut_674.mask = 64'h00ffffff7fffffff;

	lut_sub lut_680 ({sk[137], n_n980, n_n983, n_n882, n_n986, x5384x}, x5388x);
	defparam lut_680.LUT_SIZE = 6;
	defparam lut_680.mask = 64'h00ffffff7fffffff;

	lut_sub lut_686 ({sk[138], n_n1001, n_n1004, x223x, x5383x, x5386x}, x5389x);
	defparam lut_686.LUT_SIZE = 6;
	defparam lut_686.mask = 64'h00ffffff7fffffff;

	lut_sub lut_692 ({sk[139], x168x, n_n953, n_n652, x195x}, x5403x);
	defparam lut_692.LUT_SIZE = 5;
	defparam lut_692.mask = 32'h0f0f7fff;

	lut_sub lut_697 ({sk[140], x97x, x125x, x303x, x5393x, x5400x}, x5404x);
	defparam lut_697.LUT_SIZE = 6;
	defparam lut_697.mask = 64'h00ffffff7fffffff;

	lut_sub lut_703 ({sk[141], x282x, x285x, x5472x, x5474x, x5475x}, x5484x);
	defparam lut_703.LUT_SIZE = 6;
	defparam lut_703.mask = 64'h00ffffff7fffffff;

	lut_sub lut_709 ({sk[142], x119x, x160x, x5524x, x5532x, x5536x}, x5539x);
	defparam lut_709.LUT_SIZE = 6;
	defparam lut_709.mask = 64'h00ffffff7fffffff;

	lut_sub lut_715 ({sk[143], x101x, x102x, x5504x, x5505x, x5507x}, x5513x);
	defparam lut_715.LUT_SIZE = 6;
	defparam lut_715.mask = 64'h00ffffff7fffffff;

	lut_sub lut_721 ({sk[144], n_n94, x5493x, n_n1130, n_n1164, x246x}, x5508x);
	defparam lut_721.LUT_SIZE = 6;
	defparam lut_721.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_726 ({sk[145], n_n1125, x1082x, x262x, n_n1163, x265x}, x5509x);
	defparam lut_726.LUT_SIZE = 6;
	defparam lut_726.mask = 64'h00ffffff7fffffff;

	lut_sub lut_732 ({sk[146], x220x, x281x, x5526x, x5528x, x5529x}, x5538x);
	defparam lut_732.LUT_SIZE = 6;
	defparam lut_732.mask = 64'h00ffffff7fffffff;

	lut_sub lut_738 ({sk[147], x5599x, x5600x, x5601x, x5602x, x5603x}, n_n514);
	defparam lut_738.LUT_SIZE = 6;
	defparam lut_738.mask = 64'h00ffffff7fffffff;

	lut_sub lut_744 ({sk[148], n_n92, x66x, x132x, n_n71, x5668x}, x5676x);
	defparam lut_744.LUT_SIZE = 6;
	defparam lut_744.mask = 64'h00ffffff55775f7f;

	lut_sub lut_748 ({sk[149], n_n58, x36x, x224x, x1384x, x670x}, x5677x);
	defparam lut_748.LUT_SIZE = 6;
	defparam lut_748.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_753 ({sk[150], n_n95, x67x, n_n1169, x5664x, x6342x}, x5680x);
	defparam lut_753.LUT_SIZE = 6;
	defparam lut_753.mask = 64'h00ffffffbfbfbfff;

	lut_sub lut_758 ({sk[151], n_n211, x120x, x139x, x5672x, x5673x}, x5682x);
	defparam lut_758.LUT_SIZE = 6;
	defparam lut_758.mask = 64'h00ffffff7fffffff;

	lut_sub lut_764 ({sk[152], x5743x, x5744x, x5746x, x6339x}, n_n308);
	defparam lut_764.LUT_SIZE = 5;
	defparam lut_764.mask = 32'h0f0fbfff;

	lut_sub lut_769 ({sk[153], n_n1091, n_n982, x268x, x5751x, x5753x}, x5773x);
	defparam lut_769.LUT_SIZE = 6;
	defparam lut_769.mask = 64'h00ffffff7fffffff;

	lut_sub lut_775 ({sk[154], n_n84, n_n83, n_n82, x6338x, x6350x}, x5774x);
	defparam lut_775.LUT_SIZE = 6;
	defparam lut_775.mask = 64'h00ffffffeeeeeeef;

	lut_sub lut_779 ({sk[155], x162x, x266x, x5763x, x6337x}, x5776x);
	defparam lut_779.LUT_SIZE = 5;
	defparam lut_779.mask = 32'h0f0fbfff;

	lut_sub lut_784 ({sk[156], x303x, x5393x, x5769x, x5770x}, x5778x);
	defparam lut_784.LUT_SIZE = 5;
	defparam lut_784.mask = 32'h0f0f7fff;

	lut_sub lut_789 ({sk[157], x5841x, x5842x, x5844x, x6334x}, n_n376);
	defparam lut_789.LUT_SIZE = 5;
	defparam lut_789.mask = 32'h0f0fbfff;

	lut_sub lut_794 ({sk[158], n_n1286, n_n1283, x158x, x159x, x5848x}, x5869x);
	defparam lut_794.LUT_SIZE = 6;
	defparam lut_794.mask = 64'h00ffffff7fffffff;

	lut_sub lut_800 ({sk[159], x335x, x340x, x5850x, x5852x, x5853x}, x5870x);
	defparam lut_800.LUT_SIZE = 6;
	defparam lut_800.mask = 64'h00ffffff7fffffff;

	lut_sub lut_806 ({sk[160], x301x, x5858x, x5859x, x5860x}, x5872x);
	defparam lut_806.LUT_SIZE = 5;
	defparam lut_806.mask = 32'h0f0f7fff;

	lut_sub lut_811 ({sk[161], x5826x, x5827x, x5854x, x5855x, x5866x}, x5874x);
	defparam lut_811.LUT_SIZE = 6;
	defparam lut_811.mask = 64'h00ffffff7fffffff;

	lut_sub lut_817 ({sk[162], x138x, x268x, x5886x, x5892x}, x5896x);
	defparam lut_817.LUT_SIZE = 5;
	defparam lut_817.mask = 32'h0f0f7fff;

	lut_sub lut_822 ({sk[163], n_n1014, x152x, n_n1018, x5889x, x5895x}, x5897x);
	defparam lut_822.LUT_SIZE = 6;
	defparam lut_822.mask = 64'h00ffffff7fffffff;

	lut_sub lut_828 ({sk[164], x168x, n_n211, x5927x}, x5934x);
	defparam lut_828.LUT_SIZE = 4;
	defparam lut_828.mask = 16'h777f;

	lut_sub lut_832 ({sk[165], x303x, x92x, x155x, x307x, x5919x}, x5935x);
	defparam lut_832.LUT_SIZE = 6;
	defparam lut_832.mask = 64'h00ffffff7fffffff;

	lut_sub lut_838 ({sk[166], x226x, x267x, x5921x, x5922x, x5924x}, x5936x);
	defparam lut_838.LUT_SIZE = 6;
	defparam lut_838.mask = 64'h00ffffff7fffffff;

	lut_sub lut_844 ({sk[167], n_n95, n_n1079, x34x, x753x, x5609x}, x5953x);
	defparam lut_844.LUT_SIZE = 6;
	defparam lut_844.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_849 ({sk[168], n_n102, n_n94, n_n63, x282x, x287x}, x5954x);
	defparam lut_849.LUT_SIZE = 6;
	defparam lut_849.mask = 64'h00ffffff7777777f;

	lut_sub lut_853 ({sk[169], n_n1030, n_n1021, x151x, x98x, x154x}, x5955x);
	defparam lut_853.LUT_SIZE = 6;
	defparam lut_853.mask = 64'h00ffffff7fffffff;

	lut_sub lut_859 ({sk[170], n_n1057, n_n1087, x280x, x5944x, x5946x}, x5956x);
	defparam lut_859.LUT_SIZE = 6;
	defparam lut_859.mask = 64'h00ffffff7fffffff;

	lut_sub lut_865 ({sk[171], x125x, n_n652, x5990x, x5991x, x6018x}, x6026x);
	defparam lut_865.LUT_SIZE = 6;
	defparam lut_865.mask = 64'h00ffffff7fffffff;

	lut_sub lut_871 ({sk[172], n_n1215, x350x, x5964x, x5975x, x5984x}, x5987x);
	defparam lut_871.LUT_SIZE = 6;
	defparam lut_871.mask = 64'h00ffffff7fffffff;

	lut_sub lut_877 ({sk[173], n_n58, x23x, x5910x, x5514x, x6360x}, x5985x);
	defparam lut_877.LUT_SIZE = 6;
	defparam lut_877.mask = 64'h00ffffffbfbfbfff;

	lut_sub lut_882 ({sk[174], x155x, x225x, x5971x, x5972x, x5974x}, x5986x);
	defparam lut_882.LUT_SIZE = 6;
	defparam lut_882.mask = 64'h00ffffff7fffffff;

	lut_sub lut_888 ({sk[175], x6009x, x6010x, x6011x, x6012x}, x6024x);
	defparam lut_888.LUT_SIZE = 5;
	defparam lut_888.mask = 32'h0f0f7fff;

	lut_sub lut_893 ({sk[176], x6013x, x6014x, x6015x, x6016x}, x6025x);
	defparam lut_893.LUT_SIZE = 5;
	defparam lut_893.mask = 32'h0f0f7fff;

	lut_sub lut_898 ({sk[177], i_3_, i_2_, i_0_}, n_n80);
	defparam lut_898.LUT_SIZE = 4;
	defparam lut_898.mask = 16'h7740;

	lut_sub lut_900 ({sk[178], i_7_, i_8_}, n_n75);
	defparam lut_900.LUT_SIZE = 3;
	defparam lut_900.mask = 8'h54;

	lut_sub lut_902 ({sk[179], i_5_, i_4_}, x341x);
	defparam lut_902.LUT_SIZE = 3;
	defparam lut_902.mask = 8'h51;

	lut_sub lut_904 ({sk[180], i_5_, i_3_, i_4_}, n_n81);
	defparam lut_904.LUT_SIZE = 4;
	defparam lut_904.mask = 16'h7701;

	lut_sub lut_906 ({sk[181], i_7_, i_6_}, n_n38);
	defparam lut_906.LUT_SIZE = 3;
	defparam lut_906.mask = 8'h52;

	lut_sub lut_908 ({sk[182], i_7_, i_8_}, n_n64);
	defparam lut_908.LUT_SIZE = 3;
	defparam lut_908.mask = 8'h51;

	lut_sub lut_910 ({sk[183], i_7_, i_8_, i_6_}, n_n58);
	defparam lut_910.LUT_SIZE = 4;
	defparam lut_910.mask = 16'h7702;

	lut_sub lut_912 ({sk[184], i_7_, i_6_}, n_n52);
	defparam lut_912.LUT_SIZE = 3;
	defparam lut_912.mask = 8'h51;

	lut_sub lut_914 ({sk[185], i_7_, i_8_, i_6_}, n_n101);
	defparam lut_914.LUT_SIZE = 4;
	defparam lut_914.mask = 16'h7704;

	lut_sub lut_916 ({sk[186], i_7_, i_8_}, n_n86);
	defparam lut_916.LUT_SIZE = 3;
	defparam lut_916.mask = 8'h58;

	lut_sub lut_918 ({sk[187], i_7_, i_8_, i_6_}, n_n93);
	defparam lut_918.LUT_SIZE = 4;
	defparam lut_918.mask = 16'h7740;

	lut_sub lut_920 ({sk[188], i_7_, i_6_}, n_n73);
	defparam lut_920.LUT_SIZE = 3;
	defparam lut_920.mask = 8'h58;

	lut_sub lut_922 ({sk[189], i_7_, i_8_, i_6_}, n_n78);
	defparam lut_922.LUT_SIZE = 4;
	defparam lut_922.mask = 16'h7780;

	lut_sub lut_924 ({sk[190], i_7_, i_8_, i_6_}, n_n91);
	defparam lut_924.LUT_SIZE = 4;
	defparam lut_924.mask = 16'h7710;

	lut_sub lut_926 ({sk[191], i_1_, i_0_}, x175x);
	defparam lut_926.LUT_SIZE = 3;
	defparam lut_926.mask = 8'h52;

	lut_sub lut_928 ({sk[192], i_5_, i_3_, i_4_, i_2_, x175x}, x76x);
	defparam lut_928.LUT_SIZE = 6;
	defparam lut_928.mask = 64'h00ffffff10000000;

	lut_sub lut_930 ({sk[193], i_7_, i_8_, i_6_, x76x}, n_n1281);
	defparam lut_930.LUT_SIZE = 5;
	defparam lut_930.mask = 32'h0f0f0100;

	lut_sub lut_932 ({sk[194], i_1_, i_2_, i_0_}, n_n100);
	defparam lut_932.LUT_SIZE = 4;
	defparam lut_932.mask = 16'h7740;

	lut_sub lut_934 ({sk[195], i_5_, i_3_, i_4_, n_n100}, x27x);
	defparam lut_934.LUT_SIZE = 5;
	defparam lut_934.mask = 32'h0f0f0400;

	lut_sub lut_936 ({sk[196], i_5_, i_3_, i_4_, n_n78, n_n100}, n_n1185);
	defparam lut_936.LUT_SIZE = 6;
	defparam lut_936.mask = 64'h00ffffff00100000;

	lut_sub lut_938 ({sk[197], i_5_, i_3_, i_4_, i_2_, x108x}, x42x);
	defparam lut_938.LUT_SIZE = 6;
	defparam lut_938.mask = 64'h00ffffff00001000;

	lut_sub lut_940 ({sk[198], i_5_, i_3_, i_4_, n_n83, n_n95}, n_n1120);
	defparam lut_940.LUT_SIZE = 6;
	defparam lut_940.mask = 64'h00ffffff00000010;

	lut_sub lut_942 ({sk[199], i_7_, i_6_, i_3_, x341x, n_n83}, x355x);
	defparam lut_942.LUT_SIZE = 6;
	defparam lut_942.mask = 64'h00ffffff01000000;

	lut_sub lut_944 ({sk[200], i_7_, i_8_, i_6_, x128x}, n_n1156);
	defparam lut_944.LUT_SIZE = 5;
	defparam lut_944.mask = 32'h0f0f0100;

	lut_sub lut_946 ({sk[201], i_5_, i_3_, i_4_, n_n85, n_n82}, n_n1021);
	defparam lut_946.LUT_SIZE = 6;
	defparam lut_946.mask = 64'h00ffffff00001000;

	lut_sub lut_948 ({sk[202], n_n100, n_n70, n_n54, n_n1134, n_n1091}, x4837x);
	defparam lut_948.LUT_SIZE = 6;
	defparam lut_948.mask = 64'h00ffffff7777777f;

	lut_sub lut_952 ({sk[203], i_1_, i_0_}, x108x);
	defparam lut_952.LUT_SIZE = 3;
	defparam lut_952.mask = 8'h51;

	lut_sub lut_954 ({sk[204], i_5_, i_3_, i_4_, i_2_, x108x}, x57x);
	defparam lut_954.LUT_SIZE = 6;
	defparam lut_954.mask = 64'h00ffffff10000000;

	lut_sub lut_956 ({sk[205], i_5_, i_3_, i_4_}, n_n92);
	defparam lut_956.LUT_SIZE = 4;
	defparam lut_956.mask = 16'h7702;

	lut_sub lut_958 ({sk[206], i_1_, i_2_, i_0_}, n_n103);
	defparam lut_958.LUT_SIZE = 4;
	defparam lut_958.mask = 16'h7702;

	lut_sub lut_960 ({sk[207], i_5_, i_3_, i_4_, i_2_, x175x}, x26x);
	defparam lut_960.LUT_SIZE = 6;
	defparam lut_960.mask = 64'h00ffffff00000010;

	lut_sub lut_962 ({sk[208], i_5_, i_3_, i_4_}, n_n84);
	defparam lut_962.LUT_SIZE = 4;
	defparam lut_962.mask = 16'h7720;

	lut_sub lut_964 ({sk[209], i_1_, i_2_, i_0_}, n_n83);
	defparam lut_964.LUT_SIZE = 4;
	defparam lut_964.mask = 16'h7710;

	lut_sub lut_966 ({sk[210], i_1_, i_2_, i_0_, n_n91}, x32x);
	defparam lut_966.LUT_SIZE = 5;
	defparam lut_966.mask = 32'h0f0f0100;

	lut_sub lut_968 ({sk[211], i_5_, i_3_, i_4_}, n_n102);
	defparam lut_968.LUT_SIZE = 4;
	defparam lut_968.mask = 16'h7710;

	lut_sub lut_970 ({sk[212], i_1_, i_2_, i_0_}, n_n94);
	defparam lut_970.LUT_SIZE = 4;
	defparam lut_970.mask = 16'h7708;

	lut_sub lut_972 ({sk[213], i_5_, i_3_, i_4_, i_2_, x175x}, x39x);
	defparam lut_972.LUT_SIZE = 6;
	defparam lut_972.mask = 64'h00ffffff00040000;

	lut_sub lut_974 ({sk[214], i_5_, i_3_, i_4_}, n_n74);
	defparam lut_974.LUT_SIZE = 4;
	defparam lut_974.mask = 16'h7740;

	lut_sub lut_976 ({sk[215], i_1_, i_2_, i_0_}, n_n97);
	defparam lut_976.LUT_SIZE = 4;
	defparam lut_976.mask = 16'h7701;

	lut_sub lut_978 ({sk[216], i_5_, i_3_, i_4_, n_n100}, x45x);
	defparam lut_978.LUT_SIZE = 5;
	defparam lut_978.mask = 32'h0f0f0004;

	lut_sub lut_980 ({sk[217], i_5_, i_3_, i_4_, i_2_, x175x}, x55x);
	defparam lut_980.LUT_SIZE = 6;
	defparam lut_980.mask = 64'h00ffffff00004000;

	lut_sub lut_982 ({sk[218], i_5_, i_4_}, x325x);
	defparam lut_982.LUT_SIZE = 3;
	defparam lut_982.mask = 8'h54;

	lut_sub lut_984 ({sk[219], i_3_, i_1_, i_2_, i_0_, x325x}, x58x);
	defparam lut_984.LUT_SIZE = 6;
	defparam lut_984.mask = 64'h00ffffff00000100;

	lut_sub lut_986 ({sk[220], i_5_, i_3_, i_4_, n_n100}, x64x);
	defparam lut_986.LUT_SIZE = 5;
	defparam lut_986.mask = 32'h0f0f1000;

	lut_sub lut_988 ({sk[221], i_1_, i_2_}, x75x);
	defparam lut_988.LUT_SIZE = 3;
	defparam lut_988.mask = 8'h54;

	lut_sub lut_990 ({sk[222], i_1_, i_2_, i_0_, n_n101, n_n74}, n_n1217);
	defparam lut_990.LUT_SIZE = 6;
	defparam lut_990.mask = 64'h00ffffff00000010;

	lut_sub lut_992 ({sk[223], i_5_, i_3_, i_4_}, n_n77);
	defparam lut_992.LUT_SIZE = 4;
	defparam lut_992.mask = 16'h7704;

	lut_sub lut_994 ({sk[224], i_7_, i_6_, n_n97, n_n1217, n_n77}, x87x);
	defparam lut_994.LUT_SIZE = 6;
	defparam lut_994.mask = 64'h00ffffff37333333;

	lut_sub lut_997 ({sk[225], i_7_, i_8_, i_6_}, n_n95);
	defparam lut_997.LUT_SIZE = 4;
	defparam lut_997.mask = 16'h7701;

	lut_sub lut_999 ({sk[226], n_n91, n_n92, n_n100, n_n95, n_n77}, x104x);
	defparam lut_999.LUT_SIZE = 6;
	defparam lut_999.mask = 64'h00ffffff00030507;

	lut_sub lut_1002 ({sk[227], i_5_, i_3_, i_4_, i_0_, x75x}, x112x);
	defparam lut_1002.LUT_SIZE = 6;
	defparam lut_1002.mask = 64'h00ffffff00000001;

	lut_sub lut_1004 ({sk[228], i_3_, i_0_}, x56x);
	defparam lut_1004.LUT_SIZE = 3;
	defparam lut_1004.mask = 8'h51;

	lut_sub lut_1006 ({sk[229], i_7_, i_8_, i_5_, i_6_, i_4_}, x318x);
	defparam lut_1006.LUT_SIZE = 6;
	defparam lut_1006.mask = 64'h00ffffff40000000;

	lut_sub lut_1008 ({sk[230], i_5_, i_3_, i_4_, i_2_, x175x}, x63x);
	defparam lut_1008.LUT_SIZE = 6;
	defparam lut_1008.mask = 64'h00ffffff00001000;

	lut_sub lut_1010 ({sk[231], i_1_, n_n101, x56x, x318x, x63x}, x113x);
	defparam lut_1010.LUT_SIZE = 6;
	defparam lut_1010.mask = 64'h00ffffff03570055;

	lut_sub lut_1013 ({sk[232], i_7_, i_8_}, n_n70);
	defparam lut_1013.LUT_SIZE = 3;
	defparam lut_1013.mask = 8'h52;

	lut_sub lut_1015 ({sk[233], i_7_, i_8_, i_4_}, x172x);
	defparam lut_1015.LUT_SIZE = 4;
	defparam lut_1015.mask = 16'h7704;

	lut_sub lut_1017 ({sk[234], i_7_, i_8_, i_6_, i_2_, x175x}, x31x);
	defparam lut_1017.LUT_SIZE = 6;
	defparam lut_1017.mask = 64'h00ffffff04000000;

	lut_sub lut_1019 ({sk[235], n_n81, n_n103, n_n74, n_n95, x31x}, x208x);
	defparam lut_1019.LUT_SIZE = 6;
	defparam lut_1019.mask = 64'h00ffffff00035557;

	lut_sub lut_1022 ({sk[236], i_7_, i_8_, i_6_, x57x, x42x}, x227x);
	defparam lut_1022.LUT_SIZE = 6;
	defparam lut_1022.mask = 64'h00ffffff00030500;

	lut_sub lut_1025 ({sk[237], i_7_, i_8_, i_6_, x42x}, x235x);
	defparam lut_1025.LUT_SIZE = 5;
	defparam lut_1025.mask = 32'h0f0f0100;

	lut_sub lut_1027 ({sk[238], i_7_, i_8_, i_6_, n_n92, n_n103}, x252x);
	defparam lut_1027.LUT_SIZE = 6;
	defparam lut_1027.mask = 64'h00ffffff01000000;

	lut_sub lut_1029 ({sk[239], i_1_, i_2_, i_0_}, n_n85);
	defparam lut_1029.LUT_SIZE = 4;
	defparam lut_1029.mask = 16'h7704;

	lut_sub lut_1031 ({sk[240], i_6_, i_3_, i_1_, i_2_, i_0_}, x311x);
	defparam lut_1031.LUT_SIZE = 6;
	defparam lut_1031.mask = 64'h00ffffff00400000;

	lut_sub lut_1033 ({sk[241], i_5_, i_3_, i_4_, i_2_, x175x}, x25x);
	defparam lut_1033.LUT_SIZE = 6;
	defparam lut_1033.mask = 64'h00ffffff00000001;

	lut_sub lut_1035 ({sk[242], i_5_, i_3_, i_4_, n_n101, n_n103}, x329x);
	defparam lut_1035.LUT_SIZE = 6;
	defparam lut_1035.mask = 64'h00ffffff00000001;

	lut_sub lut_1037 ({sk[243], i_5_, i_6_, i_4_}, n_n54);
	defparam lut_1037.LUT_SIZE = 4;
	defparam lut_1037.mask = 16'h7708;

	lut_sub lut_1039 ({sk[244], i_7_, i_8_, i_5_, i_6_, i_4_}, x337x);
	defparam lut_1039.LUT_SIZE = 6;
	defparam lut_1039.mask = 64'h00ffffff00080000;

	lut_sub lut_1041 ({sk[245], i_5_, i_3_, i_4_, n_n1036, x107x}, x201x);
	defparam lut_1041.LUT_SIZE = 6;
	defparam lut_1041.mask = 64'h00ffffff37333333;

	lut_sub lut_1044 ({sk[246], i_3_, n_n58, n_n83, n_n95, x110x}, x164x);
	defparam lut_1044.LUT_SIZE = 6;
	defparam lut_1044.mask = 64'h00ffffff010f0000;

	lut_sub lut_1047 ({sk[247], i_7_, i_8_, i_6_, x34x, n_n1040}, x4887x);
	defparam lut_1047.LUT_SIZE = 6;
	defparam lut_1047.mask = 64'h00ffffff55555557;

	lut_sub lut_1050 ({sk[248], i_6_, n_n91, x110x, n_n67, x249x}, x4888x);
	defparam lut_1050.LUT_SIZE = 6;
	defparam lut_1050.mask = 64'h00ffffff55555557;

	lut_sub lut_1053 ({sk[249], i_7_, i_6_, x22x, x324x, x327x}, x4889x);
	defparam lut_1053.LUT_SIZE = 6;
	defparam lut_1053.mask = 64'h00ffffff11111f11;

	lut_sub lut_1056 ({sk[250], x201x, x164x, x4887x, x4888x, x4889x}, x4899x);
	defparam lut_1056.LUT_SIZE = 6;
	defparam lut_1056.mask = 64'h00ffffff7fffffff;

	lut_sub lut_1062 ({sk[251], i_5_, n_n93, n_n83, n_n1046, x288x}, x4891x);
	defparam lut_1062.LUT_SIZE = 6;
	defparam lut_1062.mask = 64'h00ffffff777f7777;

	lut_sub lut_1066 ({sk[252], i_8_, n_n58, x53x, n_n1052, x70x}, x4892x);
	defparam lut_1066.LUT_SIZE = 6;
	defparam lut_1066.mask = 64'h00ffffff777f333f;

	lut_sub lut_1070 ({sk[253], n_n82, x237x, n_n1013, x4885x, x6348x}, x4898x);
	defparam lut_1070.LUT_SIZE = 6;
	defparam lut_1070.mask = 64'h00ffffffbfbfbfff;

	lut_sub lut_1075 ({sk[254], i_2_, n_n75, x108x, n_n76, x146x}, x298x);
	defparam lut_1075.LUT_SIZE = 6;
	defparam lut_1075.mask = 64'h00ffffff55575555;

	lut_sub lut_1078 ({sk[255], n_n80, n_n70, n_n973, n_n71, n_n975}, x292x);
	defparam lut_1078.LUT_SIZE = 6;
	defparam lut_1078.mask = 64'h00ffffff5f5f5f7f;

	lut_sub lut_1082 ({sk[256], n_n78, x64x, n_n95, x29x, x1557x}, n_n882);
	defparam lut_1082.LUT_SIZE = 6;
	defparam lut_1082.mask = 64'h00ffffff555f777f;

	lut_sub lut_1086 ({sk[257], i_7_, i_0_, n_n80, n_n77, n_n943}, x4910x);
	defparam lut_1086.LUT_SIZE = 6;
	defparam lut_1086.mask = 64'h00ffffff55555575;

	lut_sub lut_1089 ({sk[258], n_n95, x41x, n_n952, n_n976, n_n986}, x4913x);
	defparam lut_1089.LUT_SIZE = 6;
	defparam lut_1089.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1094 ({sk[259], x42x, n_n95, n_n984, n_n1006, n_n978}, x4914x);
	defparam lut_1094.LUT_SIZE = 6;
	defparam lut_1094.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1099 ({sk[260], n_n982, n_n967, x204x, x202x, x203x}, x4917x);
	defparam lut_1099.LUT_SIZE = 6;
	defparam lut_1099.mask = 64'h00ffffff7fffffff;

	lut_sub lut_1105 ({sk[261], i_3_, i_4_}, x54x);
	defparam lut_1105.LUT_SIZE = 3;
	defparam lut_1105.mask = 8'h54;

	lut_sub lut_1107 ({sk[262], i_7_, i_8_, i_6_}, n_n82);
	defparam lut_1107.LUT_SIZE = 4;
	defparam lut_1107.mask = 16'h7708;

	lut_sub lut_1109 ({sk[263], i_1_, i_2_, i_0_}, n_n90);
	defparam lut_1109.LUT_SIZE = 4;
	defparam lut_1109.mask = 16'h7720;

	lut_sub lut_1111 ({sk[264], i_5_, i_3_, i_4_, n_n95, n_n90}, n_n1172);
	defparam lut_1111.LUT_SIZE = 6;
	defparam lut_1111.mask = 64'h00ffffff00000001;

	lut_sub lut_1113 ({sk[265], i_5_, i_3_, i_4_, n_n78, n_n97}, n_n1078);
	defparam lut_1113.LUT_SIZE = 6;
	defparam lut_1113.mask = 64'h00ffffff10000000;

	lut_sub lut_1115 ({sk[266], i_3_, i_2_, i_0_}, x245x);
	defparam lut_1115.LUT_SIZE = 4;
	defparam lut_1115.mask = 16'h7701;

	lut_sub lut_1117 ({sk[267], i_7_, i_8_, i_5_, i_6_, i_4_}, x38x);
	defparam lut_1117.LUT_SIZE = 6;
	defparam lut_1117.mask = 64'h00ffffff00000008;

	lut_sub lut_1119 ({sk[268], i_5_, i_3_, i_4_, i_0_, x75x}, x43x);
	defparam lut_1119.LUT_SIZE = 6;
	defparam lut_1119.mask = 64'h00ffffff04000000;

	lut_sub lut_1121 ({sk[269], i_5_, i_3_, i_4_, n_n78, n_n90}, n_n1279);
	defparam lut_1121.LUT_SIZE = 6;
	defparam lut_1121.mask = 64'h00ffffff01000000;

	lut_sub lut_1123 ({sk[270], i_7_, i_8_, i_6_, x29x, x23x}, x61x);
	defparam lut_1123.LUT_SIZE = 6;
	defparam lut_1123.mask = 64'h00ffffff00350000;

	lut_sub lut_1126 ({sk[271], i_3_, x341x, n_n94, n_n95, x239x}, x139x);
	defparam lut_1126.LUT_SIZE = 6;
	defparam lut_1126.mask = 64'h00ffffff11111113;

	lut_sub lut_1129 ({sk[272], i_1_, n_n78, x52x, x30x, x339x}, x118x);
	defparam lut_1129.LUT_SIZE = 6;
	defparam lut_1129.mask = 64'h00ffffff000f111f;

	lut_sub lut_1132 ({sk[273], n_n78, n_n91, x39x, x55x, x22x}, x6352x);
	defparam lut_1132.LUT_SIZE = 6;
	defparam lut_1132.mask = 64'h00fffffffff08880;

	lut_sub lut_1137 ({sk[274], x61x, x139x, x118x, x6352x}, n_n137);
	defparam lut_1137.LUT_SIZE = 5;
	defparam lut_1137.mask = 32'h0f0fbfff;

	lut_sub lut_1142 ({sk[275], i_8_, i_6_}, x111x);
	defparam lut_1142.LUT_SIZE = 3;
	defparam lut_1142.mask = 8'h52;

	lut_sub lut_1144 ({sk[276], i_5_, i_3_, i_4_, n_n100}, x41x);
	defparam lut_1144.LUT_SIZE = 5;
	defparam lut_1144.mask = 32'h0f0f0100;

	lut_sub lut_1146 ({sk[277], i_7_, i_8_, i_6_, x25x, x21x}, x4927x);
	defparam lut_1146.LUT_SIZE = 6;
	defparam lut_1146.mask = 64'h00ffffff30000500;

	lut_sub lut_1149 ({sk[278], i_5_, i_3_, i_4_, n_n91, n_n85}, x340x);
	defparam lut_1149.LUT_SIZE = 6;
	defparam lut_1149.mask = 64'h00ffffff00000010;

	lut_sub lut_1151 ({sk[279], n_n93, n_n102, x175x, x354x, x62x}, x4934x);
	defparam lut_1151.LUT_SIZE = 6;
	defparam lut_1151.mask = 64'h00ffffff1111111f;

	lut_sub lut_1154 ({sk[280], i_4_, n_n75, x311x, x340x, x4934x}, x4936x);
	defparam lut_1154.LUT_SIZE = 6;
	defparam lut_1154.mask = 64'h00ffffff7777777f;

	lut_sub lut_1158 ({sk[281], i_5_, i_3_, i_4_, n_n58, n_n90}, n_n1153);
	defparam lut_1158.LUT_SIZE = 6;
	defparam lut_1158.mask = 64'h00ffffff00010000;

	lut_sub lut_1160 ({sk[282], i_5_, i_3_, i_4_, i_2_, x108x}, x44x);
	defparam lut_1160.LUT_SIZE = 6;
	defparam lut_1160.mask = 64'h00ffffff00400000;

	lut_sub lut_1162 ({sk[283], i_7_, i_8_, n_n92, n_n85, n_n87}, x4938x);
	defparam lut_1162.LUT_SIZE = 6;
	defparam lut_1162.mask = 64'h00ffffff00110300;

	lut_sub lut_1165 ({sk[284], n_n58, n_n101, x57x, x25x, x350x}, x304x);
	defparam lut_1165.LUT_SIZE = 6;
	defparam lut_1165.mask = 64'h00ffffff555f777f;

	lut_sub lut_1169 ({sk[285], i_7_, i_8_, x44x, x4938x, x304x}, x4943x);
	defparam lut_1169.LUT_SIZE = 6;
	defparam lut_1169.mask = 64'h00ffffff7f777777;

	lut_sub lut_1173 ({sk[286], i_5_, i_3_, i_4_, n_n95, n_n90}, n_n1297);
	defparam lut_1173.LUT_SIZE = 6;
	defparam lut_1173.mask = 64'h00ffffff00001000;

	lut_sub lut_1175 ({sk[287], i_7_, i_8_, i_6_, n_n102, n_n90}, n_n1324);
	defparam lut_1175.LUT_SIZE = 6;
	defparam lut_1175.mask = 64'h00ffffff01000000;

	lut_sub lut_1177 ({sk[288], i_5_, i_3_, i_4_, n_n91, n_n100}, n_n1092);
	defparam lut_1177.LUT_SIZE = 6;
	defparam lut_1177.mask = 64'h00ffffff00100000;

	lut_sub lut_1179 ({sk[289], i_1_, i_2_, i_0_, n_n102, n_n95}, n_n1103);
	defparam lut_1179.LUT_SIZE = 6;
	defparam lut_1179.mask = 64'h00ffffff00010000;

	lut_sub lut_1181 ({sk[290], i_7_, i_5_, i_6_, x54x, n_n90}, x319x);
	defparam lut_1181.LUT_SIZE = 6;
	defparam lut_1181.mask = 64'h00ffffff00100000;

	lut_sub lut_1183 ({sk[291], i_7_, i_8_, i_6_, n_n84, n_n85}, n_n1130);
	defparam lut_1183.LUT_SIZE = 6;
	defparam lut_1183.mask = 64'h00ffffff00000010;

	lut_sub lut_1185 ({sk[292], i_5_, i_6_, i_3_}, x354x);
	defparam lut_1185.LUT_SIZE = 4;
	defparam lut_1185.mask = 16'h7740;

	lut_sub lut_1187 ({sk[293], i_7_, i_8_, i_1_, i_2_, i_0_}, x4944x);
	defparam lut_1187.LUT_SIZE = 6;
	defparam lut_1187.mask = 64'h00ffffff00000800;

	lut_sub lut_1189 ({sk[294], n_n1103, x319x, n_n1130, x354x, x4944x}, x4950x);
	defparam lut_1189.LUT_SIZE = 6;
	defparam lut_1189.mask = 64'h00ffffff1fffffff;

	lut_sub lut_1194 ({sk[295], i_5_, i_3_, i_4_, n_n58, n_n94}, n_n1105);
	defparam lut_1194.LUT_SIZE = 6;
	defparam lut_1194.mask = 64'h00ffffff00000001;

	lut_sub lut_1196 ({sk[296], i_5_, i_3_, i_4_, n_n93, n_n90}, n_n1108);
	defparam lut_1196.LUT_SIZE = 6;
	defparam lut_1196.mask = 64'h00ffffff00000001;

	lut_sub lut_1198 ({sk[297], i_7_, i_8_, n_n84, n_n83, n_n1100}, x94x);
	defparam lut_1198.LUT_SIZE = 6;
	defparam lut_1198.mask = 64'h00ffffff55555557;

	lut_sub lut_1201 ({sk[298], n_n63, x44x, n_n1105, n_n1108, x94x}, x4951x);
	defparam lut_1201.LUT_SIZE = 6;
	defparam lut_1201.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1206 ({sk[299], i_5_, i_1_, i_2_, i_0_, x54x}, x19x);
	defparam lut_1206.LUT_SIZE = 6;
	defparam lut_1206.mask = 64'h00ffffff00000004;

	lut_sub lut_1208 ({sk[300], i_5_, i_3_, i_4_, i_2_, x108x}, x29x);
	defparam lut_1208.LUT_SIZE = 6;
	defparam lut_1208.mask = 64'h00ffffff00010000;

	lut_sub lut_1210 ({sk[301], i_1_, i_2_, i_0_, n_n38, n_n70}, x37x);
	defparam lut_1210.LUT_SIZE = 6;
	defparam lut_1210.mask = 64'h00ffffff00001000;

	lut_sub lut_1212 ({sk[302], n_n81, n_n91, n_n100, n_n83, n_n74}, x105x);
	defparam lut_1212.LUT_SIZE = 6;
	defparam lut_1212.mask = 64'h00ffffff0011001f;

	lut_sub lut_1215 ({sk[303], i_5_, i_4_}, x109x);
	defparam lut_1215.LUT_SIZE = 3;
	defparam lut_1215.mask = 8'h52;

	lut_sub lut_1217 ({sk[304], i_6_, i_3_, i_4_}, x127x);
	defparam lut_1217.LUT_SIZE = 4;
	defparam lut_1217.mask = 16'h7704;

	lut_sub lut_1219 ({sk[305], i_5_, i_3_, i_4_, n_n97, n_n63}, n_n1082);
	defparam lut_1219.LUT_SIZE = 6;
	defparam lut_1219.mask = 64'h00ffffff01000000;

	lut_sub lut_1221 ({sk[306], i_5_, i_4_}, x110x);
	defparam lut_1221.LUT_SIZE = 3;
	defparam lut_1221.mask = 8'h58;

	lut_sub lut_1223 ({sk[307], i_7_, i_6_, i_3_, n_n83, x110x}, x1487x);
	defparam lut_1223.LUT_SIZE = 6;
	defparam lut_1223.mask = 64'h00ffffff10000000;

	lut_sub lut_1225 ({sk[308], n_n75, n_n38, n_n84, x55x, n_n90}, x207x);
	defparam lut_1225.LUT_SIZE = 6;
	defparam lut_1225.mask = 64'h00ffffff00053337;

	lut_sub lut_1228 ({sk[309], i_7_, i_8_, i_3_, n_n103, x109x}, x1483x);
	defparam lut_1228.LUT_SIZE = 6;
	defparam lut_1228.mask = 64'h00ffffff00100000;

	lut_sub lut_1230 ({sk[310], i_7_, i_8_, i_3_, n_n85, x325x}, x1484x);
	defparam lut_1230.LUT_SIZE = 6;
	defparam lut_1230.mask = 64'h00ffffff00000100;

	lut_sub lut_1232 ({sk[311], i_3_, i_1_, i_0_}, n_n67);
	defparam lut_1232.LUT_SIZE = 4;
	defparam lut_1232.mask = 16'h7740;

	lut_sub lut_1234 ({sk[312], i_7_, i_6_, i_2_, n_n102, x175x}, x1479x);
	defparam lut_1234.LUT_SIZE = 6;
	defparam lut_1234.mask = 64'h00ffffff00000100;

	lut_sub lut_1236 ({sk[313], i_1_, i_2_, i_0_, x35x}, x1480x);
	defparam lut_1236.LUT_SIZE = 5;
	defparam lut_1236.mask = 32'h0f0f0100;

	lut_sub lut_1238 ({sk[314], i_7_, i_8_, i_6_, n_n103, n_n77}, x251x);
	defparam lut_1238.LUT_SIZE = 6;
	defparam lut_1238.mask = 64'h00ffffff00100000;

	lut_sub lut_1240 ({sk[315], i_7_, i_8_, i_6_, n_n81, n_n100}, n_n1079);
	defparam lut_1240.LUT_SIZE = 6;
	defparam lut_1240.mask = 64'h00ffffff01000000;

	lut_sub lut_1242 ({sk[316], i_5_, i_3_, i_4_, n_n1079, x31x}, x254x);
	defparam lut_1242.LUT_SIZE = 6;
	defparam lut_1242.mask = 64'h00ffffff73333333;

	lut_sub lut_1245 ({sk[317], i_5_, i_3_, i_4_, n_n101, n_n97}, x321x);
	defparam lut_1245.LUT_SIZE = 6;
	defparam lut_1245.mask = 64'h00ffffff01000000;

	lut_sub lut_1247 ({sk[318], i_7_, i_8_, i_1_, i_2_, i_0_}, x328x);
	defparam lut_1247.LUT_SIZE = 6;
	defparam lut_1247.mask = 64'h00ffffff00000001;

	lut_sub lut_1249 ({sk[319], i_7_, i_8_, i_6_, n_n92, n_n90}, n_n1259);
	defparam lut_1249.LUT_SIZE = 6;
	defparam lut_1249.mask = 64'h00ffffff00100000;

	lut_sub lut_1251 ({sk[320], i_5_, i_3_, i_4_, n_n100}, x239x);
	defparam lut_1251.LUT_SIZE = 5;
	defparam lut_1251.mask = 32'h0f0f0040;

	lut_sub lut_1253 ({sk[321], i_7_, i_8_, i_6_, x239x}, n_n1204);
	defparam lut_1253.LUT_SIZE = 5;
	defparam lut_1253.mask = 32'h0f0f0001;

	lut_sub lut_1255 ({sk[322], i_3_, i_1_, i_0_}, x351x);
	defparam lut_1255.LUT_SIZE = 4;
	defparam lut_1255.mask = 16'h7780;

	lut_sub lut_1257 ({sk[323], i_5_, i_3_, i_4_, i_0_, x75x}, x21x);
	defparam lut_1257.LUT_SIZE = 6;
	defparam lut_1257.mask = 64'h00ffffff10000000;

	lut_sub lut_1259 ({sk[324], i_3_, n_n58, n_n94, x109x, n_n1085}, x256x);
	defparam lut_1259.LUT_SIZE = 6;
	defparam lut_1259.mask = 64'h00ffffff55575555;

	lut_sub lut_1262 ({sk[325], i_6_, n_n86, x43x, n_n1040, x114x}, x299x);
	defparam lut_1262.LUT_SIZE = 6;
	defparam lut_1262.mask = 64'h00ffffff7777777f;

	lut_sub lut_1266 ({sk[326], n_n102, n_n1095, x20x, n_n1088, n_n1181}, x5006x);
	defparam lut_1266.LUT_SIZE = 6;
	defparam lut_1266.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_1271 ({sk[327], i_5_, i_3_, i_4_, x32x, n_n1160}, x190x);
	defparam lut_1271.LUT_SIZE = 6;
	defparam lut_1271.mask = 64'h00ffffff55755555;

	lut_sub lut_1274 ({sk[328], i_7_, i_8_, i_6_, x63x, n_n1146}, x265x);
	defparam lut_1274.LUT_SIZE = 6;
	defparam lut_1274.mask = 64'h00ffffff75555555;

	lut_sub lut_1277 ({sk[329], n_n58, x64x, n_n1132, x335x, x1440x}, x5003x);
	defparam lut_1277.LUT_SIZE = 6;
	defparam lut_1277.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1282 ({sk[330], x337x, n_n1172, n_n1022, x322x, n_n1128}, x5004x);
	defparam lut_1282.LUT_SIZE = 6;
	defparam lut_1282.mask = 64'h00ffffff5fff7fff;

	lut_sub lut_1287 ({sk[331], n_n58, n_n1036, x44x, n_n1060, n_n1164}, x5005x);
	defparam lut_1287.LUT_SIZE = 6;
	defparam lut_1287.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_1292 ({sk[332], i_4_, i_1_, i_2_, i_0_, x28x}, x135x);
	defparam lut_1292.LUT_SIZE = 6;
	defparam lut_1292.mask = 64'h00ffffffc400c000;

	lut_sub lut_1295 ({sk[333], i_5_, i_3_, i_4_, n_n101, n_n85}, n_n949);
	defparam lut_1295.LUT_SIZE = 6;
	defparam lut_1295.mask = 64'h00ffffff00100000;

	lut_sub lut_1297 ({sk[334], i_7_, i_8_, i_6_, x49x, n_n941}, x97x);
	defparam lut_1297.LUT_SIZE = 6;
	defparam lut_1297.mask = 64'h00ffffff57555555;

	lut_sub lut_1300 ({sk[335], i_7_, i_8_, i_6_, x52x, n_n951}, x204x);
	defparam lut_1300.LUT_SIZE = 6;
	defparam lut_1300.mask = 64'h00ffffff55555557;

	lut_sub lut_1303 ({sk[336], x25x, n_n82, n_n1021, x249x, n_n978}, x5025x);
	defparam lut_1303.LUT_SIZE = 6;
	defparam lut_1303.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1308 ({sk[337], i_0_, n_n78, x75x, x42x, x5012x}, x195x);
	defparam lut_1308.LUT_SIZE = 6;
	defparam lut_1308.mask = 64'h00ffffff05370033;

	lut_sub lut_1311 ({sk[338], i_3_, x341x, n_n78, n_n100, n_n1018}, x151x);
	defparam lut_1311.LUT_SIZE = 6;
	defparam lut_1311.mask = 64'h00ffffff55555557;

	lut_sub lut_1314 ({sk[339], n_n103, n_n74, n_n82, x79x, n_n975}, x5021x);
	defparam lut_1314.LUT_SIZE = 6;
	defparam lut_1314.mask = 64'h00ffffff7777777f;

	lut_sub lut_1318 ({sk[340], n_n78, x29x, n_n967, n_n969, x1557x}, x5023x);
	defparam lut_1318.LUT_SIZE = 6;
	defparam lut_1318.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1323 ({sk[341], n_n95, x41x, x128x, x44x, n_n1004}, x5024x);
	defparam lut_1323.LUT_SIZE = 6;
	defparam lut_1323.mask = 64'h00ffffff55557fff;

	lut_sub lut_1328 ({sk[342], i_5_, i_3_, i_4_, i_2_, x108x}, x34x);
	defparam lut_1328.LUT_SIZE = 6;
	defparam lut_1328.mask = 64'h00ffffff40000000;

	lut_sub lut_1330 ({sk[343], i_5_, i_3_, i_4_, i_2_, x108x}, x23x);
	defparam lut_1330.LUT_SIZE = 6;
	defparam lut_1330.mask = 64'h00ffffff00000001;

	lut_sub lut_1332 ({sk[344], i_5_, i_3_, i_4_, n_n58, n_n90}, n_n1188);
	defparam lut_1332.LUT_SIZE = 6;
	defparam lut_1332.mask = 64'h00ffffff00000001;

	lut_sub lut_1334 ({sk[345], i_6_, n_n86, n_n74, n_n97, n_n1188}, x88x);
	defparam lut_1334.LUT_SIZE = 6;
	defparam lut_1334.mask = 64'h00ffffff55555557;

	lut_sub lut_1337 ({sk[346], i_5_, i_3_, i_4_, n_n100, n_n82}, x346x);
	defparam lut_1337.LUT_SIZE = 6;
	defparam lut_1337.mask = 64'h00ffffff01000000;

	lut_sub lut_1339 ({sk[347], i_5_, i_3_, i_4_, n_n103, n_n82}, x1413x);
	defparam lut_1339.LUT_SIZE = 6;
	defparam lut_1339.mask = 64'h00ffffff00000010;

	lut_sub lut_1341 ({sk[348], i_7_, i_8_, i_6_, n_n81, n_n97}, x1414x);
	defparam lut_1341.LUT_SIZE = 6;
	defparam lut_1341.mask = 64'h00ffffff00100000;

	lut_sub lut_1343 ({sk[349], i_5_, i_3_, i_4_, n_n101, n_n103}, x343x);
	defparam lut_1343.LUT_SIZE = 6;
	defparam lut_1343.mask = 64'h00ffffff00000010;

	lut_sub lut_1345 ({sk[350], i_7_, i_8_, i_6_, x34x}, x1518x);
	defparam lut_1345.LUT_SIZE = 5;
	defparam lut_1345.mask = 32'h0f0f0040;

	lut_sub lut_1347 ({sk[351], i_5_, i_3_, i_4_, n_n58, n_n100}, x1519x);
	defparam lut_1347.LUT_SIZE = 6;
	defparam lut_1347.mask = 64'h00ffffff00000100;

	lut_sub lut_1349 ({sk[352], i_3_, x38x, x108x, x1518x, x1519x}, x231x);
	defparam lut_1349.LUT_SIZE = 6;
	defparam lut_1349.mask = 64'h00ffffff777f7777;

	lut_sub lut_1353 ({sk[353], i_7_, i_8_, i_6_, n_n84, n_n94}, n_n1193);
	defparam lut_1353.LUT_SIZE = 6;
	defparam lut_1353.mask = 64'h00ffffff00000010;

	lut_sub lut_1355 ({sk[354], n_n58, n_n78, n_n100, n_n84, n_n94}, x255x);
	defparam lut_1355.LUT_SIZE = 6;
	defparam lut_1355.mask = 64'h00ffffff00031113;

	lut_sub lut_1358 ({sk[355], i_5_, i_3_, i_4_, i_2_, x108x}, x46x);
	defparam lut_1358.LUT_SIZE = 6;
	defparam lut_1358.mask = 64'h00ffffff00000040;

	lut_sub lut_1360 ({sk[356], i_7_, i_8_, i_6_, x46x, x41x}, x5031x);
	defparam lut_1360.LUT_SIZE = 6;
	defparam lut_1360.mask = 64'h00ffffff05000003;

	lut_sub lut_1363 ({sk[357], i_7_, i_8_, i_6_, x21x, x5031x}, x301x);
	defparam lut_1363.LUT_SIZE = 6;
	defparam lut_1363.mask = 64'h00ffffff55575555;

	lut_sub lut_1366 ({sk[358], i_5_, i_3_, i_4_, i_2_, x108x}, x53x);
	defparam lut_1366.LUT_SIZE = 6;
	defparam lut_1366.mask = 64'h00ffffff00040000;

	lut_sub lut_1368 ({sk[359], i_7_, i_8_, i_6_, n_n102, n_n85}, n_n1022);
	defparam lut_1368.LUT_SIZE = 6;
	defparam lut_1368.mask = 64'h00ffffff00000010;

	lut_sub lut_1370 ({sk[360], i_7_, i_8_, i_6_, n_n100, n_n74}, n_n1134);
	defparam lut_1370.LUT_SIZE = 6;
	defparam lut_1370.mask = 64'h00ffffff00000010;

	lut_sub lut_1372 ({sk[361], i_5_, i_3_, i_4_, n_n78, n_n94}, n_n1039);
	defparam lut_1372.LUT_SIZE = 6;
	defparam lut_1372.mask = 64'h00ffffff00010000;

	lut_sub lut_1374 ({sk[362], i_7_, i_8_, i_5_, i_6_, i_4_}, x78x);
	defparam lut_1374.LUT_SIZE = 6;
	defparam lut_1374.mask = 64'h00ffffff00000004;

	lut_sub lut_1376 ({sk[363], i_5_, i_6_, i_4_}, n_n87);
	defparam lut_1376.LUT_SIZE = 4;
	defparam lut_1376.mask = 16'h7704;

	lut_sub lut_1378 ({sk[364], i_3_, i_2_, i_0_, n_n64, n_n87}, n_n1091);
	defparam lut_1378.LUT_SIZE = 6;
	defparam lut_1378.mask = 64'h00ffffff00000100;

	lut_sub lut_1380 ({sk[365], n_n58, x25x, n_n1153, n_n1267, x342x}, x5060x);
	defparam lut_1380.LUT_SIZE = 6;
	defparam lut_1380.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1385 ({sk[366], n_n95, x67x, n_n1216, n_n1146, n_n1164}, x5061x);
	defparam lut_1385.LUT_SIZE = 6;
	defparam lut_1385.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1390 ({sk[367], n_n101, n_n92, n_n103, n_n1170, x5056x}, x5062x);
	defparam lut_1390.LUT_SIZE = 6;
	defparam lut_1390.mask = 64'h00ffffff7777777f;

	lut_sub lut_1394 ({sk[368], x87x, x61x, x224x, x1384x}, x5063x);
	defparam lut_1394.LUT_SIZE = 5;
	defparam lut_1394.mask = 32'h0f0f7fff;

	lut_sub lut_1399 ({sk[369], x206x, x225x, x5059x}, x5064x);
	defparam lut_1399.LUT_SIZE = 4;
	defparam lut_1399.mask = 16'h777f;

	lut_sub lut_1403 ({sk[370], x42x, n_n95, n_n983, n_n999, x249x}, x5076x);
	defparam lut_1403.LUT_SIZE = 6;
	defparam lut_1403.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1408 ({sk[371], n_n951, n_n954, n_n952, x147x, x202x}, x5077x);
	defparam lut_1408.LUT_SIZE = 6;
	defparam lut_1408.mask = 64'h00ffffff7fffffff;

	lut_sub lut_1414 ({sk[372], x294x, x146x, n_n1001, n_n1010, n_n978}, x5078x);
	defparam lut_1414.LUT_SIZE = 6;
	defparam lut_1414.mask = 64'h00ffffff7fffffff;

	lut_sub lut_1420 ({sk[373], x97x, n_n939, n_n981, x272x, x151x}, x5079x);
	defparam lut_1420.LUT_SIZE = 6;
	defparam lut_1420.mask = 64'h00ffffff7fffffff;

	lut_sub lut_1426 ({sk[374], i_3_, i_2_, i_0_}, x322x);
	defparam lut_1426.LUT_SIZE = 4;
	defparam lut_1426.mask = 16'h7720;

	lut_sub lut_1428 ({sk[375], i_7_, i_8_, i_6_, x109x, x322x}, n_n1093);
	defparam lut_1428.LUT_SIZE = 6;
	defparam lut_1428.mask = 64'h00ffffff00100000;

	lut_sub lut_1430 ({sk[376], i_1_, i_2_, i_0_, n_n74, n_n63}, n_n1052);
	defparam lut_1430.LUT_SIZE = 6;
	defparam lut_1430.mask = 64'h00ffffff00001000;

	lut_sub lut_1432 ({sk[377], i_5_, i_3_, i_4_, n_n91, n_n90}, n_n1331);
	defparam lut_1432.LUT_SIZE = 6;
	defparam lut_1432.mask = 64'h00ffffff01000000;

	lut_sub lut_1434 ({sk[378], i_5_, i_6_, i_4_}, n_n40);
	defparam lut_1434.LUT_SIZE = 4;
	defparam lut_1434.mask = 16'h7740;

	lut_sub lut_1436 ({sk[379], i_3_, n_n75, n_n38, x109x, n_n40}, x35x);
	defparam lut_1436.LUT_SIZE = 6;
	defparam lut_1436.mask = 64'h00ffffff03570055;

	lut_sub lut_1439 ({sk[380], i_5_, i_3_, i_4_, n_n94, n_n82}, x1359x);
	defparam lut_1439.LUT_SIZE = 6;
	defparam lut_1439.mask = 64'h00ffffff01000000;

	lut_sub lut_1441 ({sk[381], i_5_, i_6_, i_4_}, n_n66);
	defparam lut_1441.LUT_SIZE = 4;
	defparam lut_1441.mask = 16'h7702;

	lut_sub lut_1443 ({sk[382], i_7_, i_8_, i_6_, i_2_, x108x}, x20x);
	defparam lut_1443.LUT_SIZE = 6;
	defparam lut_1443.mask = 64'h00ffffff04000000;

	lut_sub lut_1445 ({sk[383], i_3_, i_1_, i_2_}, x353x);
	defparam lut_1445.LUT_SIZE = 4;
	defparam lut_1445.mask = 16'h7740;

	lut_sub lut_1447 ({sk[384], n_n86, n_n77, n_n66, x20x, x353x}, x117x);
	defparam lut_1447.LUT_SIZE = 6;
	defparam lut_1447.mask = 64'h00ffffff00330537;

	lut_sub lut_1450 ({sk[385], i_1_, i_2_, i_0_, n_n58, n_n74}, n_n1058);
	defparam lut_1450.LUT_SIZE = 6;
	defparam lut_1450.mask = 64'h00ffffff00001000;

	lut_sub lut_1452 ({sk[386], i_7_, i_6_, n_n103, n_n84, n_n1058}, x133x);
	defparam lut_1452.LUT_SIZE = 6;
	defparam lut_1452.mask = 64'h00ffffff55555755;

	lut_sub lut_1455 ({sk[387], i_7_, i_8_, i_6_, n_n74, n_n90}, n_n1032);
	defparam lut_1455.LUT_SIZE = 6;
	defparam lut_1455.mask = 64'h00ffffff01000000;

	lut_sub lut_1457 ({sk[388], i_5_, i_3_, i_4_, n_n85, n_n95}, n_n1040);
	defparam lut_1457.LUT_SIZE = 6;
	defparam lut_1457.mask = 64'h00ffffff00001000;

	lut_sub lut_1459 ({sk[389], i_7_, i_8_, i_6_, x43x, n_n1040}, x148x);
	defparam lut_1459.LUT_SIZE = 6;
	defparam lut_1459.mask = 64'h00ffffff57555555;

	lut_sub lut_1462 ({sk[390], i_7_, i_6_}, x173x);
	defparam lut_1462.LUT_SIZE = 3;
	defparam lut_1462.mask = 8'h54;

	lut_sub lut_1464 ({sk[391], i_7_, i_8_, i_6_}, x177x);
	defparam lut_1464.LUT_SIZE = 4;
	defparam lut_1464.mask = 16'h7714;

	lut_sub lut_1467 ({sk[392], i_5_, i_3_, i_4_, n_n94, n_n82}, x323x);
	defparam lut_1467.LUT_SIZE = 6;
	defparam lut_1467.mask = 64'h00ffffff10000000;

	lut_sub lut_1469 ({sk[393], i_5_, i_3_, i_4_, n_n100, n_n95}, x1352x);
	defparam lut_1469.LUT_SIZE = 6;
	defparam lut_1469.mask = 64'h00ffffff00100000;

	lut_sub lut_1471 ({sk[394], i_1_, i_2_, i_0_, n_n91, n_n74}, n_n1036);
	defparam lut_1471.LUT_SIZE = 6;
	defparam lut_1471.mask = 64'h00ffffff00000010;

	lut_sub lut_1473 ({sk[395], i_1_, i_2_, i_0_, n_n101}, x107x);
	defparam lut_1473.LUT_SIZE = 5;
	defparam lut_1473.mask = 32'h0f0f0010;

	lut_sub lut_1475 ({sk[396], n_n58, n_n91, n_n103, n_n77, n_n90}, x233x);
	defparam lut_1475.LUT_SIZE = 6;
	defparam lut_1475.mask = 64'h00ffffff00031313;

	lut_sub lut_1479 ({sk[397], i_5_, i_3_, i_4_, n_n94, n_n63}, n_n1085);
	defparam lut_1479.LUT_SIZE = 6;
	defparam lut_1479.mask = 64'h00ffffff00010000;

	lut_sub lut_1481 ({sk[398], i_7_, i_6_, n_n97, n_n1078, n_n77}, x5083x);
	defparam lut_1481.LUT_SIZE = 6;
	defparam lut_1481.mask = 64'h00ffffff33333337;

	lut_sub lut_1484 ({sk[399], i_7_, i_6_, i_3_, n_n100, x110x}, x1348x);
	defparam lut_1484.LUT_SIZE = 6;
	defparam lut_1484.mask = 64'h00ffffff10000000;

	lut_sub lut_1486 ({sk[400], n_n101, n_n74, n_n90, x5083x, x1348x}, x257x);
	defparam lut_1486.LUT_SIZE = 6;
	defparam lut_1486.mask = 64'h00ffffff7777777f;

	lut_sub lut_1490 ({sk[401], i_5_, i_1_, i_2_, i_0_, x54x}, x237x);
	defparam lut_1490.LUT_SIZE = 6;
	defparam lut_1490.mask = 64'h00ffffff01000000;

	lut_sub lut_1492 ({sk[402], i_7_, i_8_, i_6_, i_3_, i_4_}, x5085x);
	defparam lut_1492.LUT_SIZE = 6;
	defparam lut_1492.mask = 64'h00ffffff00000100;

	lut_sub lut_1494 ({sk[403], i_2_, n_n82, x175x, x237x, x5085x}, x271x);
	defparam lut_1494.LUT_SIZE = 6;
	defparam lut_1494.mask = 64'h00ffffff05370033;

	lut_sub lut_1497 ({sk[404], n_n84, n_n83, n_n82, n_n983, n_n986}, x296x);
	defparam lut_1497.LUT_SIZE = 6;
	defparam lut_1497.mask = 64'h00ffffff7777777f;

	lut_sub lut_1501 ({sk[405], n_n95, x41x, n_n949, n_n969, n_n966}, x5121x);
	defparam lut_1501.LUT_SIZE = 6;
	defparam lut_1501.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1506 ({sk[406], x271x, n_n944, x145x, x146x, n_n939}, x5123x);
	defparam lut_1506.LUT_SIZE = 6;
	defparam lut_1506.mask = 64'h00ffffff7fffffff;

	lut_sub lut_1512 ({sk[407], x189x, n_n958, x270x, x272x, x5114x}, x5124x);
	defparam lut_1512.LUT_SIZE = 6;
	defparam lut_1512.mask = 64'h00ffffff7fffffff;

	lut_sub lut_1518 ({sk[408], i_3_, i_1_, i_2_, i_0_, x325x}, x52x);
	defparam lut_1518.LUT_SIZE = 6;
	defparam lut_1518.mask = 64'h00ffffff00000004;

	lut_sub lut_1520 ({sk[409], n_n93, x57x, n_n63, x83x, n_n1177}, x306x);
	defparam lut_1520.LUT_SIZE = 6;
	defparam lut_1520.mask = 64'h00ffffff575757ff;

	lut_sub lut_1524 ({sk[410], i_6_, n_n86, x257x, n_n1158, x65x}, x5135x);
	defparam lut_1524.LUT_SIZE = 6;
	defparam lut_1524.mask = 64'h00ffffff3f3f3f7f;

	lut_sub lut_1528 ({sk[411], i_3_, n_n52, x39x, x110x, x31x}, x141x);
	defparam lut_1528.LUT_SIZE = 6;
	defparam lut_1528.mask = 64'h00ffffff111f000f;

	lut_sub lut_1531 ({sk[412], i_0_, n_n102, x75x, n_n95, n_n1095}, x279x);
	defparam lut_1531.LUT_SIZE = 6;
	defparam lut_1531.mask = 64'h00ffffff55555557;

	lut_sub lut_1534 ({sk[413], i_8_, i_6_, n_n81, n_n85, x133x}, x5131x);
	defparam lut_1534.LUT_SIZE = 6;
	defparam lut_1534.mask = 64'h00ffffff55555755;

	lut_sub lut_1537 ({sk[414], n_n91, n_n100, n_n84, n_n1153, x267x}, x5133x);
	defparam lut_1537.LUT_SIZE = 6;
	defparam lut_1537.mask = 64'h00ffffff7777777f;

	lut_sub lut_1541 ({sk[415], n_n74, n_n1082, n_n1120, n_n1052, x107x}, x5134x);
	defparam lut_1541.LUT_SIZE = 6;
	defparam lut_1541.mask = 64'h00ffffff3fff7fff;

	lut_sub lut_1546 ({sk[416], i_5_, i_3_, i_4_, i_2_, x175x}, x67x);
	defparam lut_1546.LUT_SIZE = 6;
	defparam lut_1546.mask = 64'h00ffffff00400000;

	lut_sub lut_1548 ({sk[417], i_5_, i_3_, i_4_, n_n95, n_n90}, n_n1330);
	defparam lut_1548.LUT_SIZE = 6;
	defparam lut_1548.mask = 64'h00ffffff00010000;

	lut_sub lut_1550 ({sk[418], i_5_, i_3_, i_4_, n_n101, n_n100}, n_n1267);
	defparam lut_1550.LUT_SIZE = 6;
	defparam lut_1550.mask = 64'h00ffffff00100000;

	lut_sub lut_1552 ({sk[419], i_5_, i_3_, i_4_, i_0_, x75x}, x36x);
	defparam lut_1552.LUT_SIZE = 6;
	defparam lut_1552.mask = 64'h00ffffff00000400;

	lut_sub lut_1554 ({sk[420], i_1_, i_2_, i_0_, n_n73, x111x}, x48x);
	defparam lut_1554.LUT_SIZE = 6;
	defparam lut_1554.mask = 64'h00ffffff00010000;

	lut_sub lut_1556 ({sk[421], i_7_, i_5_, i_3_, i_4_, i_0_}, x72x);
	defparam lut_1556.LUT_SIZE = 6;
	defparam lut_1556.mask = 64'h00ffffff80008080;

	lut_sub lut_1559 ({sk[422], i_1_, i_2_, i_0_, n_n101, n_n84}, x1291x);
	defparam lut_1559.LUT_SIZE = 6;
	defparam lut_1559.mask = 64'h00ffffff00000010;

	lut_sub lut_1561 ({sk[423], i_5_, i_3_, i_4_, n_n93, n_n85}, x1292x);
	defparam lut_1561.LUT_SIZE = 6;
	defparam lut_1561.mask = 64'h00ffffff00000010;

	lut_sub lut_1563 ({sk[424], i_2_, i_0_}, x327x);
	defparam lut_1563.LUT_SIZE = 3;
	defparam lut_1563.mask = 8'h51;

	lut_sub lut_1565 ({sk[425], i_3_, n_n93, x38x, x19x, x327x}, x123x);
	defparam lut_1565.LUT_SIZE = 6;
	defparam lut_1565.mask = 64'h00ffffff05370033;

	lut_sub lut_1568 ({sk[426], n_n93, x76x, n_n84, n_n63, n_n90}, x183x);
	defparam lut_1568.LUT_SIZE = 6;
	defparam lut_1568.mask = 64'h00ffffff00330537;

	lut_sub lut_1571 ({sk[427], i_5_, i_3_, i_4_, n_n78, n_n97}, x1285x);
	defparam lut_1571.LUT_SIZE = 6;
	defparam lut_1571.mask = 64'h00ffffff01000000;

	lut_sub lut_1573 ({sk[428], i_5_, i_3_, i_4_, n_n78, n_n100}, x348x);
	defparam lut_1573.LUT_SIZE = 6;
	defparam lut_1573.mask = 64'h00ffffff00000100;

	lut_sub lut_1575 ({sk[429], i_5_, i_3_, i_4_, i_2_, x175x}, x128x);
	defparam lut_1575.LUT_SIZE = 6;
	defparam lut_1575.mask = 64'h00ffffff40000000;

	lut_sub lut_1577 ({sk[430], i_7_, i_8_, i_6_, x348x, x128x}, x186x);
	defparam lut_1577.LUT_SIZE = 6;
	defparam lut_1577.mask = 64'h00ffffff33333373;

	lut_sub lut_1580 ({sk[431], i_2_, n_n101, n_n84, x108x, x78x}, x206x);
	defparam lut_1580.LUT_SIZE = 6;
	defparam lut_1580.mask = 64'h00ffffff11110003;

	lut_sub lut_1583 ({sk[432], i_5_, i_6_, i_3_}, n_n76);
	defparam lut_1583.LUT_SIZE = 4;
	defparam lut_1583.mask = 16'h7704;

	lut_sub lut_1585 ({sk[433], i_7_, i_8_, i_6_, x239x}, n_n1215);
	defparam lut_1585.LUT_SIZE = 5;
	defparam lut_1585.mask = 32'h0f0f0004;

	lut_sub lut_1587 ({sk[434], i_7_, i_6_, i_2_, n_n77, x175x}, x342x);
	defparam lut_1587.LUT_SIZE = 6;
	defparam lut_1587.mask = 64'h00ffffff10000000;

	lut_sub lut_1589 ({sk[435], i_7_, i_6_, n_n1082, x21x, x52x}, x5176x);
	defparam lut_1589.LUT_SIZE = 6;
	defparam lut_1589.mask = 64'h00ffffff3f0f5f0f;

	lut_sub lut_1593 ({sk[436], x48x, n_n1216, n_n1088, n_n1181, x194x}, x5181x);
	defparam lut_1593.LUT_SIZE = 6;
	defparam lut_1593.mask = 64'h00ffffff3fff7fff;

	lut_sub lut_1598 ({sk[437], i_7_, i_6_, x34x, n_n1215, x190x}, x5178x);
	defparam lut_1598.LUT_SIZE = 6;
	defparam lut_1598.mask = 64'h00ffffff7777777f;

	lut_sub lut_1602 ({sk[438], n_n100, n_n1204, x78x, n_n1128, n_n1184}, x5179x);
	defparam lut_1602.LUT_SIZE = 6;
	defparam lut_1602.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_1607 ({sk[439], n_n91, x63x, n_n1132, n_n1130, x335x}, x5180x);
	defparam lut_1607.LUT_SIZE = 6;
	defparam lut_1607.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1612 ({sk[440], n_n101, x42x, n_n95, n_n942, x52x}, x125x);
	defparam lut_1612.LUT_SIZE = 6;
	defparam lut_1612.mask = 64'h00ffffff333f777f;

	lut_sub lut_1616 ({sk[441], i_2_, x38x, x108x, n_n973, n_n975}, x5193x);
	defparam lut_1616.LUT_SIZE = 6;
	defparam lut_1616.mask = 64'h00ffffff777f7777;

	lut_sub lut_1620 ({sk[442], n_n95, x52x, x128x, n_n986, n_n1042}, x5198x);
	defparam lut_1620.LUT_SIZE = 6;
	defparam lut_1620.mask = 64'h00ffffff77777fff;

	lut_sub lut_1625 ({sk[443], n_n91, x29x, x189x, n_n958, n_n1060}, x5196x);
	defparam lut_1625.LUT_SIZE = 6;
	defparam lut_1625.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1630 ({sk[444], x64x, n_n95, n_n980, n_n999, n_n1004}, x5197x);
	defparam lut_1630.LUT_SIZE = 6;
	defparam lut_1630.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1635 ({sk[445], n_n967, n_n966, x147x, x195x, x274x}, x5200x);
	defparam lut_1635.LUT_SIZE = 6;
	defparam lut_1635.mask = 64'h00ffffff7fffffff;

	lut_sub lut_1641 ({sk[446], i_7_, i_8_, i_1_, i_2_, i_0_}, x62x);
	defparam lut_1641.LUT_SIZE = 6;
	defparam lut_1641.mask = 64'h00ffffff10000000;

	lut_sub lut_1643 ({sk[447], i_6_, n_n91, x34x, x110x, x62x}, x185x);
	defparam lut_1643.LUT_SIZE = 6;
	defparam lut_1643.mask = 64'h00ffffff111f000f;

	lut_sub lut_1646 ({sk[448], i_5_, i_3_, i_4_, n_n78, n_n90}, x352x);
	defparam lut_1646.LUT_SIZE = 6;
	defparam lut_1646.mask = 64'h00ffffff00001000;

	lut_sub lut_1648 ({sk[449], i_1_, i_2_, i_0_, n_n101, n_n74}, n_n1074);
	defparam lut_1648.LUT_SIZE = 6;
	defparam lut_1648.mask = 64'h00ffffff00001000;

	lut_sub lut_1650 ({sk[450], i_5_, i_3_, i_4_, n_n78, n_n90}, n_n1294);
	defparam lut_1650.LUT_SIZE = 6;
	defparam lut_1650.mask = 64'h00ffffff00100000;

	lut_sub lut_1652 ({sk[451], i_5_, i_3_, i_4_, n_n101, n_n90}, n_n1109);
	defparam lut_1652.LUT_SIZE = 6;
	defparam lut_1652.mask = 64'h00ffffff01000000;

	lut_sub lut_1654 ({sk[452], i_5_, i_3_, i_4_, n_n93, n_n90}, n_n1132);
	defparam lut_1654.LUT_SIZE = 6;
	defparam lut_1654.mask = 64'h00ffffff00001000;

	lut_sub lut_1656 ({sk[453], i_6_, i_3_}, x28x);
	defparam lut_1656.LUT_SIZE = 3;
	defparam lut_1656.mask = 8'h58;

	lut_sub lut_1658 ({sk[454], i_6_, i_3_, i_4_}, x131x);
	defparam lut_1658.LUT_SIZE = 4;
	defparam lut_1658.mask = 16'h7780;

	lut_sub lut_1660 ({sk[455], i_5_, i_6_, i_3_, i_4_}, x5012x);
	defparam lut_1660.LUT_SIZE = 5;
	defparam lut_1660.mask = 32'h0f0f0800;

	lut_sub lut_1662 ({sk[456], i_5_, i_3_, i_4_, n_n101, n_n90}, n_n1312);
	defparam lut_1662.LUT_SIZE = 6;
	defparam lut_1662.mask = 64'h00ffffff00001000;

	lut_sub lut_1664 ({sk[457], i_1_, i_2_, i_0_, n_n101, n_n77}, x326x);
	defparam lut_1664.LUT_SIZE = 6;
	defparam lut_1664.mask = 64'h00ffffff00001000;

	lut_sub lut_1666 ({sk[458], i_5_, i_3_, i_4_, n_n91, n_n90}, n_n1169);
	defparam lut_1666.LUT_SIZE = 6;
	defparam lut_1666.mask = 64'h00ffffff00010000;

	lut_sub lut_1668 ({sk[459], i_5_, i_3_, i_4_, n_n91, n_n94}, n_n942);
	defparam lut_1668.LUT_SIZE = 6;
	defparam lut_1668.mask = 64'h00ffffff00000010;

	lut_sub lut_1670 ({sk[460], i_5_, i_3_, i_4_, n_n82, n_n90}, n_n1057);
	defparam lut_1670.LUT_SIZE = 6;
	defparam lut_1670.mask = 64'h00ffffff00000001;

	lut_sub lut_1672 ({sk[461], i_5_, i_3_, i_4_, n_n78, n_n90}, n_n1125);
	defparam lut_1672.LUT_SIZE = 6;
	defparam lut_1672.mask = 64'h00ffffff00000001;

	lut_sub lut_1674 ({sk[462], i_5_, i_3_, i_4_, n_n78, n_n94}, n_n1128);
	defparam lut_1674.LUT_SIZE = 6;
	defparam lut_1674.mask = 64'h00ffffff00100000;

	lut_sub lut_1676 ({sk[463], i_7_, i_6_, i_3_, n_n94, x109x}, x333x);
	defparam lut_1676.LUT_SIZE = 6;
	defparam lut_1676.mask = 64'h00ffffff00000001;

	lut_sub lut_1678 ({sk[464], i_5_, i_3_, i_4_, n_n58, n_n94}, n_n1286);
	defparam lut_1678.LUT_SIZE = 6;
	defparam lut_1678.mask = 64'h00ffffff00000010;

	lut_sub lut_1680 ({sk[465], i_7_, i_6_, n_n74, n_n90, n_n1286}, x278x);
	defparam lut_1680.LUT_SIZE = 6;
	defparam lut_1680.mask = 64'h00ffffff55555755;

	lut_sub lut_1683 ({sk[466], i_5_, i_3_, i_4_, n_n63, n_n90}, n_n1047);
	defparam lut_1683.LUT_SIZE = 6;
	defparam lut_1683.mask = 64'h00ffffff00000001;

	lut_sub lut_1685 ({sk[467], i_7_, i_8_, i_6_, n_n92, n_n94}, n_n1042);
	defparam lut_1685.LUT_SIZE = 6;
	defparam lut_1685.mask = 64'h00ffffff01000000;

	lut_sub lut_1687 ({sk[468], i_1_, i_2_, i_0_}, n_n937);
	defparam lut_1687.LUT_SIZE = 4;
	defparam lut_1687.mask = 16'h7780;

	lut_sub lut_1689 ({sk[469], i_5_, i_6_, i_4_, x351x, n_n937}, x189x);
	defparam lut_1689.LUT_SIZE = 6;
	defparam lut_1689.mask = 64'h00ffffff75555555;

	lut_sub lut_1692 ({sk[470], i_5_, i_3_, i_4_, n_n93, n_n94}, n_n941);
	defparam lut_1692.LUT_SIZE = 6;
	defparam lut_1692.mask = 64'h00ffffff00001000;

	lut_sub lut_1694 ({sk[471], i_5_, i_3_, i_4_, n_n94, n_n63}, n_n1087);
	defparam lut_1694.LUT_SIZE = 6;
	defparam lut_1694.mask = 64'h00ffffff00000001;

	lut_sub lut_1696 ({sk[472], n_n101, n_n83, n_n102, x1359x, x217x}, x5273x);
	defparam lut_1696.LUT_SIZE = 6;
	defparam lut_1696.mask = 64'h00ffffff7777777f;

	lut_sub lut_1700 ({sk[473], i_2_, x56x, x318x, n_n1294, x290x}, x5274x);
	defparam lut_1700.LUT_SIZE = 6;
	defparam lut_1700.mask = 64'h00ffffff777f7777;

	lut_sub lut_1704 ({sk[474], i_6_, n_n86, x27x, x4938x, x6349x}, x5306x);
	defparam lut_1704.LUT_SIZE = 6;
	defparam lut_1704.mask = 64'h00ffffffbbbbbbbf;

	lut_sub lut_1708 ({sk[475], x227x, n_n77, x207x, x61x, x20x}, x5307x);
	defparam lut_1708.LUT_SIZE = 6;
	defparam lut_1708.mask = 64'h00ffffff3f7fffff;

	lut_sub lut_1713 ({sk[476], n_n101, x55x, x323x, x1352x, x1143x}, x5298x);
	defparam lut_1713.LUT_SIZE = 6;
	defparam lut_1713.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1718 ({sk[477], x352x, n_n1176, x5283x, x6346x}, x5309x);
	defparam lut_1718.LUT_SIZE = 5;
	defparam lut_1718.mask = 32'h0f0fbfff;

	lut_sub lut_1723 ({sk[478], x333x, x332x, x5288x, x5289x, x5290x}, x5310x);
	defparam lut_1723.LUT_SIZE = 6;
	defparam lut_1723.mask = 64'h00ffffff7fffffff;

	lut_sub lut_1729 ({sk[479], x71x, x118x, x5291x, x5292x, x5305x}, x6345x);
	defparam lut_1729.LUT_SIZE = 6;
	defparam lut_1729.mask = 64'h00ffffff80000000;

	lut_sub lut_1731 ({sk[480], i_7_, i_8_, i_5_, i_6_, i_4_}, x234x);
	defparam lut_1731.LUT_SIZE = 6;
	defparam lut_1731.mask = 64'h00ffffff00002000;

	lut_sub lut_1733 ({sk[481], i_1_, i_2_, i_0_, n_n95, n_n77}, n_n958);
	defparam lut_1733.LUT_SIZE = 6;
	defparam lut_1733.mask = 64'h00ffffff00000100;

	lut_sub lut_1735 ({sk[482], i_7_, i_8_, i_5_, i_6_, i_4_}, x320x);
	defparam lut_1735.LUT_SIZE = 6;
	defparam lut_1735.mask = 64'h00ffffff00000200;

	lut_sub lut_1737 ({sk[483], i_1_, i_2_, i_0_, n_n74, n_n82}, n_n973);
	defparam lut_1737.LUT_SIZE = 6;
	defparam lut_1737.mask = 64'h00ffffff00000010;

	lut_sub lut_1739 ({sk[484], i_5_, i_3_, i_4_, n_n91, n_n94}, n_n989);
	defparam lut_1739.LUT_SIZE = 6;
	defparam lut_1739.mask = 64'h00ffffff00000001;

	lut_sub lut_1741 ({sk[485], i_5_, i_3_, i_4_, n_n91, n_n97}, n_n944);
	defparam lut_1741.LUT_SIZE = 6;
	defparam lut_1741.mask = 64'h00ffffff00010000;

	lut_sub lut_1743 ({sk[486], i_7_, i_8_, i_6_, n_n81, n_n83}, n_n982);
	defparam lut_1743.LUT_SIZE = 6;
	defparam lut_1743.mask = 64'h00ffffff01000000;

	lut_sub lut_1745 ({sk[487], i_7_, i_8_, i_6_, n_n100, n_n77}, n_n967);
	defparam lut_1745.LUT_SIZE = 6;
	defparam lut_1745.mask = 64'h00ffffff01000000;

	lut_sub lut_1747 ({sk[488], i_5_, i_6_, i_4_, n_n70, n_n90}, n_n1121);
	defparam lut_1747.LUT_SIZE = 6;
	defparam lut_1747.mask = 64'h00ffffff00000001;

	lut_sub lut_1749 ({sk[489], i_3_, i_1_, i_2_}, n_n53);
	defparam lut_1749.LUT_SIZE = 4;
	defparam lut_1749.mask = 16'h7710;

	lut_sub lut_1751 ({sk[490], i_5_, i_6_, i_4_, n_n80}, x1588x);
	defparam lut_1751.LUT_SIZE = 5;
	defparam lut_1751.mask = 32'h0f0f1000;

	lut_sub lut_1753 ({sk[491], i_1_, i_2_}, x330x);
	defparam lut_1753.LUT_SIZE = 3;
	defparam lut_1753.mask = 8'h52;

	lut_sub lut_1755 ({sk[492], i_5_, i_3_, n_n73, x1588x, x330x}, x70x);
	defparam lut_1755.LUT_SIZE = 6;
	defparam lut_1755.mask = 64'h00ffffff37333333;

	lut_sub lut_1758 ({sk[493], i_5_, i_3_, i_4_, i_2_, x108x}, x83x);
	defparam lut_1758.LUT_SIZE = 6;
	defparam lut_1758.mask = 64'h00ffffff00000010;

	lut_sub lut_1760 ({sk[494], i_8_, i_6_, i_3_, n_n94, x109x}, x1082x);
	defparam lut_1760.LUT_SIZE = 6;
	defparam lut_1760.mask = 64'h00ffffff10000000;

	lut_sub lut_1762 ({sk[495], i_8_, i_6_, x55x, n_n1125}, x90x);
	defparam lut_1762.LUT_SIZE = 5;
	defparam lut_1762.mask = 32'h0f0f7555;

	lut_sub lut_1765 ({sk[496], i_1_, i_2_, i_0_, n_n78, n_n74}, n_n962);
	defparam lut_1765.LUT_SIZE = 6;
	defparam lut_1765.mask = 64'h00ffffff00010000;

	lut_sub lut_1767 ({sk[497], n_n64, n_n52, x41x, x128x, n_n962}, x168x);
	defparam lut_1767.LUT_SIZE = 6;
	defparam lut_1767.mask = 64'h00ffffff5555557f;

	lut_sub lut_1771 ({sk[498], i_5_, i_6_, i_4_}, x5338x);
	defparam lut_1771.LUT_SIZE = 4;
	defparam lut_1771.mask = 16'h7701;

	lut_sub lut_1773 ({sk[499], i_7_, i_8_, i_5_, i_6_, i_4_}, x324x);
	defparam lut_1773.LUT_SIZE = 6;
	defparam lut_1773.mask = 64'h00ffffff00000080;

	lut_sub lut_1775 ({sk[500], n_n75, n_n85, x5338x, x324x, n_n67}, x215x);
	defparam lut_1775.LUT_SIZE = 6;
	defparam lut_1775.mask = 64'h00ffffff1111111f;

	lut_sub lut_1778 ({sk[501], i_7_, i_8_, i_6_, x341x, n_n100}, x236x);
	defparam lut_1778.LUT_SIZE = 6;
	defparam lut_1778.mask = 64'h00ffffff00000010;

	lut_sub lut_1780 ({sk[502], i_7_, i_8_, i_6_, x54x, n_n90}, n_n1118);
	defparam lut_1780.LUT_SIZE = 6;
	defparam lut_1780.mask = 64'h00ffffff00010000;

	lut_sub lut_1782 ({sk[503], i_7_, i_8_, n_n84, n_n94, n_n1118}, x262x);
	defparam lut_1782.LUT_SIZE = 6;
	defparam lut_1782.mask = 64'h00ffffff55555755;

	lut_sub lut_1785 ({sk[504], i_7_, i_8_, i_6_, x25x, x237x}, x275x);
	defparam lut_1785.LUT_SIZE = 6;
	defparam lut_1785.mask = 64'h00ffffff03030005;

	lut_sub lut_1788 ({sk[505], i_5_, i_3_, i_4_, n_n85, n_n82}, n_n952);
	defparam lut_1788.LUT_SIZE = 6;
	defparam lut_1788.mask = 64'h00ffffff00000001;

	lut_sub lut_1790 ({sk[506], i_3_, x341x, n_n78, n_n94, n_n952}, x145x);
	defparam lut_1790.LUT_SIZE = 6;
	defparam lut_1790.mask = 64'h00ffffff55555557;

	lut_sub lut_1793 ({sk[507], i_5_, i_3_, i_4_, n_n83, n_n82}, n_n951);
	defparam lut_1793.LUT_SIZE = 6;
	defparam lut_1793.mask = 64'h00ffffff00000010;

	lut_sub lut_1795 ({sk[508], i_5_, i_3_, i_4_, n_n91, n_n97}, n_n959);
	defparam lut_1795.LUT_SIZE = 6;
	defparam lut_1795.mask = 64'h00ffffff00100000;

	lut_sub lut_1797 ({sk[509], i_3_, n_n91, n_n100, x109x, n_n959}, x146x);
	defparam lut_1797.LUT_SIZE = 6;
	defparam lut_1797.mask = 64'h00ffffff55555557;

	lut_sub lut_1800 ({sk[510], i_5_, i_3_, i_4_, n_n83, n_n82}, n_n980);
	defparam lut_1800.LUT_SIZE = 6;
	defparam lut_1800.mask = 64'h00ffffff00100000;

	lut_sub lut_1802 ({sk[511], i_5_, i_3_, i_4_, n_n100, n_n95}, n_n983);
	defparam lut_1802.LUT_SIZE = 6;
	defparam lut_1802.mask = 64'h00ffffff10000000;

	lut_sub lut_1804 ({sk[512], i_5_, i_3_, i_4_, n_n94, n_n63}, n_n986);
	defparam lut_1804.LUT_SIZE = 6;
	defparam lut_1804.mask = 64'h00ffffff00000010;

	lut_sub lut_1806 ({sk[513], i_3_, n_n64, x292x, x238x, x313x}, x5384x);
	defparam lut_1806.LUT_SIZE = 6;
	defparam lut_1806.mask = 64'h00ffffff0f3f5f7f;

	lut_sub lut_1810 ({sk[514], i_7_, i_8_, i_6_, x57x}, n_n1001);
	defparam lut_1810.LUT_SIZE = 5;
	defparam lut_1810.mask = 32'h0f0f0400;

	lut_sub lut_1812 ({sk[515], i_5_, i_3_, i_4_, n_n91, n_n97}, n_n1004);
	defparam lut_1812.LUT_SIZE = 6;
	defparam lut_1812.mask = 64'h00ffffff01000000;

	lut_sub lut_1814 ({sk[516], i_7_, i_8_, n_n969, n_n66, n_n67}, x223x);
	defparam lut_1814.LUT_SIZE = 6;
	defparam lut_1814.mask = 64'h00ffffff0f0f1f0f;

	lut_sub lut_1817 ({sk[517], n_n82, x237x, n_n976, n_n987, n_n994}, x5383x);
	defparam lut_1817.LUT_SIZE = 6;
	defparam lut_1817.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1822 ({sk[518], x275x, x59x, x163x, x200x}, x5386x);
	defparam lut_1822.LUT_SIZE = 5;
	defparam lut_1822.mask = 32'h0f0f7fff;

	lut_sub lut_1827 ({sk[519], i_7_, i_8_, i_6_, n_n80, x110x}, n_n953);
	defparam lut_1827.LUT_SIZE = 6;
	defparam lut_1827.mask = 64'h00ffffff10000000;

	lut_sub lut_1829 ({sk[520], n_n103, n_n102, n_n97, n_n95, n_n949}, n_n652);
	defparam lut_1829.LUT_SIZE = 6;
	defparam lut_1829.mask = 64'h00ffffff55575577;

	lut_sub lut_1833 ({sk[521], n_n73, x53x, n_n967, n_n966, x1017x}, x303x);
	defparam lut_1833.LUT_SIZE = 6;
	defparam lut_1833.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1838 ({sk[522], n_n951, n_n954, n_n952, x5392x}, x5393x);
	defparam lut_1838.LUT_SIZE = 5;
	defparam lut_1838.mask = 32'h0f0f7fff;

	lut_sub lut_1843 ({sk[523], n_n91, n_n102, n_n97, n_n939, x5399x}, x5400x);
	defparam lut_1843.LUT_SIZE = 6;
	defparam lut_1843.mask = 64'h00ffffff7777777f;

	lut_sub lut_1847 ({sk[524], i_8_, i_6_, i_3_, n_n94, x110x}, n_n1045);
	defparam lut_1847.LUT_SIZE = 6;
	defparam lut_1847.mask = 64'h00ffffff00000100;

	lut_sub lut_1849 ({sk[525], i_5_, i_3_, i_4_, n_n91, n_n85}, n_n1043);
	defparam lut_1849.LUT_SIZE = 6;
	defparam lut_1849.mask = 64'h00ffffff00010000;

	lut_sub lut_1851 ({sk[526], x27x, n_n74, n_n82, x31x, x1153x}, x290x);
	defparam lut_1851.LUT_SIZE = 6;
	defparam lut_1851.mask = 64'h00ffffff55775f7f;

	lut_sub lut_1855 ({sk[527], n_n93, n_n103, n_n74, x352x, x5407x}, x309x);
	defparam lut_1855.LUT_SIZE = 6;
	defparam lut_1855.mask = 64'h00ffffff7777777f;

	lut_sub lut_1859 ({sk[528], n_n92, x32x, n_n77, x31x, x289x}, x5417x);
	defparam lut_1859.LUT_SIZE = 6;
	defparam lut_1859.mask = 64'h00ffffff575757ff;

	lut_sub lut_1863 ({sk[529], x290x, x309x, x5417x}, x5421x);
	defparam lut_1863.LUT_SIZE = 4;
	defparam lut_1863.mask = 16'h777f;

	lut_sub lut_1867 ({sk[530], i_7_, i_8_, i_6_, x27x, x208x}, x5413x);
	defparam lut_1867.LUT_SIZE = 6;
	defparam lut_1867.mask = 64'h00ffffff57555555;

	lut_sub lut_1870 ({sk[531], n_n58, x26x, x32x, n_n102, x210x}, x5414x);
	defparam lut_1870.LUT_SIZE = 6;
	defparam lut_1870.mask = 64'h00ffffff575757ff;

	lut_sub lut_1874 ({sk[532], n_n101, n_n1281, x346x, x63x, x248x}, x5415x);
	defparam lut_1874.LUT_SIZE = 6;
	defparam lut_1874.mask = 64'h00ffffff5fff7fff;

	lut_sub lut_1879 ({sk[533], n_n64, n_n52, x57x, x326x, x5411x}, x5416x);
	defparam lut_1879.LUT_SIZE = 6;
	defparam lut_1879.mask = 64'h00ffffff7777777f;

	lut_sub lut_1883 ({sk[534], x5413x, x5414x, x5415x, x5416x}, x5422x);
	defparam lut_1883.LUT_SIZE = 5;
	defparam lut_1883.mask = 32'h0f0f7fff;

	lut_sub lut_1888 ({sk[535], i_3_, i_1_, i_2_, i_0_, x110x}, x22x);
	defparam lut_1888.LUT_SIZE = 6;
	defparam lut_1888.mask = 64'h00ffffff00000004;

	lut_sub lut_1890 ({sk[536], i_5_, n_n91, x67x, x28x, x62x}, x158x);
	defparam lut_1890.LUT_SIZE = 6;
	defparam lut_1890.mask = 64'h00ffffff000f111f;

	lut_sub lut_1893 ({sk[537], n_n58, n_n78, x23x, x33x, x5429x}, x5436x);
	defparam lut_1893.LUT_SIZE = 6;
	defparam lut_1893.mask = 64'h00ffffff555f777f;

	lut_sub lut_1897 ({sk[538], n_n101, x22x, x158x, x304x, x5436x}, x5440x);
	defparam lut_1897.LUT_SIZE = 6;
	defparam lut_1897.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_1902 ({sk[539], n_n38, n_n70, x34x, x119x, x1519x}, x5432x);
	defparam lut_1902.LUT_SIZE = 6;
	defparam lut_1902.mask = 64'h00ffffff7777777f;

	lut_sub lut_1906 ({sk[540], i_6_, n_n86, x57x, n_n1177, x122x}, x5433x);
	defparam lut_1906.LUT_SIZE = 6;
	defparam lut_1906.mask = 64'h00ffffff7777777f;

	lut_sub lut_1910 ({sk[541], n_n93, x26x, x329x, n_n1176, x22x}, x5434x);
	defparam lut_1910.LUT_SIZE = 6;
	defparam lut_1910.mask = 64'h00ffffff3f3f7fff;

	lut_sub lut_1915 ({sk[542], n_n78, x55x, x22x, x332x, n_n1170}, x5435x);
	defparam lut_1915.LUT_SIZE = 6;
	defparam lut_1915.mask = 64'h00ffffff77777fff;

	lut_sub lut_1920 ({sk[543], x5432x, x5433x, x5434x, x5435x}, x5441x);
	defparam lut_1920.LUT_SIZE = 5;
	defparam lut_1920.mask = 32'h0f0f7fff;

	lut_sub lut_1925 ({sk[544], i_5_, i_3_, i_4_, n_n83, n_n82}, n_n1030);
	defparam lut_1925.LUT_SIZE = 6;
	defparam lut_1925.mask = 64'h00ffffff00000001;

	lut_sub lut_1927 ({sk[545], i_7_, i_8_, i_1_, i_2_, i_0_}, x66x);
	defparam lut_1927.LUT_SIZE = 6;
	defparam lut_1927.mask = 64'h00ffffff00000002;

	lut_sub lut_1929 ({sk[546], i_6_, i_3_, i_4_}, x5442x);
	defparam lut_1929.LUT_SIZE = 4;
	defparam lut_1929.mask = 16'h7702;

	lut_sub lut_1931 ({sk[547], i_7_, i_8_, i_6_, x109x, x322x}, n_n1101);
	defparam lut_1931.LUT_SIZE = 6;
	defparam lut_1931.mask = 64'h00ffffff00001000;

	lut_sub lut_1933 ({sk[548], i_5_, n_n101, x58x, n_n82, x353x}, x6359x);
	defparam lut_1933.LUT_SIZE = 6;
	defparam lut_1933.mask = 64'h00fffffffca8fcfc;

	lut_sub lut_1940 ({sk[549], n_n63, n_n1128, x44x, n_n1156, x6359x}, x5450x);
	defparam lut_1940.LUT_SIZE = 6;
	defparam lut_1940.mask = 64'h00ffffffbbffbfff;

	lut_sub lut_1945 ({sk[550], i_7_, i_8_, i_0_, n_n71, x30x}, n_n1059);
	defparam lut_1945.LUT_SIZE = 6;
	defparam lut_1945.mask = 64'h00ffffff01000000;

	lut_sub lut_1947 ({sk[551], i_8_, i_1_, x56x, n_n40, n_n1060}, x156x);
	defparam lut_1947.LUT_SIZE = 6;
	defparam lut_1947.mask = 64'h00ffffff55555755;

	lut_sub lut_1950 ({sk[552], n_n38, n_n1058, n_n1059, x22x, x156x}, x5454x);
	defparam lut_1950.LUT_SIZE = 6;
	defparam lut_1950.mask = 64'h00ffffff5fff7fff;

	lut_sub lut_1955 ({sk[553], i_7_, i_8_, i_6_, x76x}, x334x);
	defparam lut_1955.LUT_SIZE = 5;
	defparam lut_1955.mask = 32'h0f0f4000;

	lut_sub lut_1957 ({sk[554], i_6_, n_n70, x110x, n_n53, x334x}, x142x);
	defparam lut_1957.LUT_SIZE = 6;
	defparam lut_1957.mask = 64'h00ffffff55575555;

	lut_sub lut_1960 ({sk[555], i_7_, i_8_, i_6_, x42x}, x944x);
	defparam lut_1960.LUT_SIZE = 5;
	defparam lut_1960.mask = 32'h0f0f0400;

	lut_sub lut_1962 ({sk[556], i_7_, i_8_, i_6_, x42x, n_n1105}, x150x);
	defparam lut_1962.LUT_SIZE = 6;
	defparam lut_1962.mask = 64'h00ffffff55755555;

	lut_sub lut_1965 ({sk[557], i_5_, i_3_, i_4_, n_n101, n_n90}, n_n1046);
	defparam lut_1965.LUT_SIZE = 6;
	defparam lut_1965.mask = 64'h00ffffff00010000;

	lut_sub lut_1967 ({sk[558], i_5_, i_3_, i_4_, n_n91, n_n103}, n_n1095);
	defparam lut_1967.LUT_SIZE = 6;
	defparam lut_1967.mask = 64'h00ffffff00000010;

	lut_sub lut_1969 ({sk[559], i_7_, i_8_, i_3_, i_1_, i_0_}, x85x);
	defparam lut_1969.LUT_SIZE = 6;
	defparam lut_1969.mask = 64'h00ffffff00400000;

	lut_sub lut_1971 ({sk[560], i_6_, x55x, n_n95, x110x, x85x}, x282x);
	defparam lut_1971.LUT_SIZE = 6;
	defparam lut_1971.mask = 64'h00ffffff000f111f;

	lut_sub lut_1974 ({sk[561], i_5_, n_n91, n_n100, x54x, n_n1074}, x285x);
	defparam lut_1974.LUT_SIZE = 6;
	defparam lut_1974.mask = 64'h00ffffff55575555;

	lut_sub lut_1977 ({sk[562], i_1_, i_2_, i_0_, n_n74, n_n63}, n_n1060);
	defparam lut_1977.LUT_SIZE = 6;
	defparam lut_1977.mask = 64'h00ffffff00000010;

	lut_sub lut_1979 ({sk[563], i_5_, i_3_, i_4_, n_n100, n_n82}, n_n1100);
	defparam lut_1979.LUT_SIZE = 6;
	defparam lut_1979.mask = 64'h00ffffff00000100;

	lut_sub lut_1981 ({sk[564], i_7_, i_8_, i_6_, i_0_, x75x}, x132x);
	defparam lut_1981.LUT_SIZE = 6;
	defparam lut_1981.mask = 64'h00ffffff01000000;

	lut_sub lut_1983 ({sk[565], i_5_, i_3_, i_4_, n_n93, n_n83}, n_n969);
	defparam lut_1983.LUT_SIZE = 6;
	defparam lut_1983.mask = 64'h00ffffff00000100;

	lut_sub lut_1985 ({sk[566], i_5_, i_3_, i_4_, n_n78, n_n94}, n_n954);
	defparam lut_1985.LUT_SIZE = 6;
	defparam lut_1985.mask = 64'h00ffffff00000001;

	lut_sub lut_1987 ({sk[567], i_8_, i_6_}, x331x);
	defparam lut_1987.LUT_SIZE = 3;
	defparam lut_1987.mask = 8'h58;

	lut_sub lut_1989 ({sk[568], i_5_, i_3_, i_4_, n_n100, x331x}, n_n939);
	defparam lut_1989.LUT_SIZE = 6;
	defparam lut_1989.mask = 64'h00ffffff10000000;

	lut_sub lut_1991 ({sk[569], i_7_, i_8_, i_1_, i_2_, i_0_}, x5068x);
	defparam lut_1991.LUT_SIZE = 6;
	defparam lut_1991.mask = 64'h00ffffff40000000;

	lut_sub lut_1993 ({sk[570], i_6_, i_3_, i_4_, n_n86, n_n100}, n_n971);
	defparam lut_1993.LUT_SIZE = 6;
	defparam lut_1993.mask = 64'h00ffffff10000000;

	lut_sub lut_1995 ({sk[571], i_8_, i_6_, i_3_, n_n94, x325x}, n_n1037);
	defparam lut_1995.LUT_SIZE = 6;
	defparam lut_1995.mask = 64'h00ffffff00010000;

	lut_sub lut_1997 ({sk[572], i_5_, i_6_, i_4_, n_n64, n_n103}, x903x);
	defparam lut_1997.LUT_SIZE = 6;
	defparam lut_1997.mask = 64'h00ffffff01000000;

	lut_sub lut_1999 ({sk[573], i_7_, i_8_, i_6_, x76x, x21x}, x5492x);
	defparam lut_1999.LUT_SIZE = 6;
	defparam lut_1999.mask = 64'h00ffffff30000005;

	lut_sub lut_2002 ({sk[574], n_n38, n_n64, x27x, n_n71, x242x}, x119x);
	defparam lut_2002.LUT_SIZE = 6;
	defparam lut_2002.mask = 64'h00ffffff0011001f;

	lut_sub lut_2005 ({sk[575], i_7_, i_8_, i_6_, x237x, x33x}, x160x);
	defparam lut_2005.LUT_SIZE = 6;
	defparam lut_2005.mask = 64'h00ffffff03000350;

	lut_sub lut_2008 ({sk[576], i_6_, n_n86, x25x, x267x, x877x}, x5524x);
	defparam lut_2008.LUT_SIZE = 6;
	defparam lut_2008.mask = 64'h00ffffff7777777f;

	lut_sub lut_2012 ({sk[577], n_n81, x32x, x278x, x159x, x5514x}, x5532x);
	defparam lut_2012.LUT_SIZE = 6;
	defparam lut_2012.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2017 ({sk[578], n_n101, x49x, x835x, x5519x, x5531x}, x5536x);
	defparam lut_2017.LUT_SIZE = 6;
	defparam lut_2017.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2022 ({sk[579], i_3_, i_1_, i_0_, n_n86, n_n87}, n_n947);
	defparam lut_2022.LUT_SIZE = 6;
	defparam lut_2022.mask = 64'h00ffffff00100000;

	lut_sub lut_2024 ({sk[580], i_7_, i_8_, i_6_, x29x, n_n947}, x162x);
	defparam lut_2024.LUT_SIZE = 6;
	defparam lut_2024.mask = 64'h00ffffff55555557;

	lut_sub lut_2027 ({sk[581], i_8_, i_6_, i_3_, i_4_, n_n97}, x829x);
	defparam lut_2027.LUT_SIZE = 6;
	defparam lut_2027.mask = 64'h00ffffff00040000;

	lut_sub lut_2029 ({sk[582], n_n92, n_n94, n_n63, n_n983, x212x}, x5550x);
	defparam lut_2029.LUT_SIZE = 6;
	defparam lut_2029.mask = 64'h00ffffff7777777f;

	lut_sub lut_2033 ({sk[583], n_n82, x237x, n_n994, n_n1013, n_n978}, x5551x);
	defparam lut_2033.LUT_SIZE = 6;
	defparam lut_2033.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2038 ({sk[584], n_n86, n_n85, n_n76, n_n882, n_n1026}, x5552x);
	defparam lut_2038.LUT_SIZE = 6;
	defparam lut_2038.mask = 64'h00ffffff7777777f;

	lut_sub lut_2042 ({sk[585], n_n987, n_n984, n_n1011, x59x, x202x}, x5553x);
	defparam lut_2042.LUT_SIZE = 6;
	defparam lut_2042.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2048 ({sk[586], n_n71, x270x, x85x, x200x, x152x}, x5554x);
	defparam lut_2048.LUT_SIZE = 6;
	defparam lut_2048.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_2053 ({sk[587], i_5_, i_6_, i_4_}, n_n71);
	defparam lut_2053.LUT_SIZE = 4;
	defparam lut_2053.mask = 16'h7720;

	lut_sub lut_2055 ({sk[588], i_3_, i_2_}, x30x);
	defparam lut_2055.LUT_SIZE = 3;
	defparam lut_2055.mask = 8'h51;

	lut_sub lut_2057 ({sk[589], i_2_, n_n70, x38x, x108x, n_n87}, x68x);
	defparam lut_2057.LUT_SIZE = 6;
	defparam lut_2057.mask = 64'h00ffffff03030011;

	lut_sub lut_2060 ({sk[590], n_n91, x54x, x108x, n_n87, x85x}, x138x);
	defparam lut_2060.LUT_SIZE = 6;
	defparam lut_2060.mask = 64'h00ffffff1111111f;

	lut_sub lut_2063 ({sk[591], i_7_, i_8_, i_6_, n_n102, n_n97}, x805x);
	defparam lut_2063.LUT_SIZE = 6;
	defparam lut_2063.mask = 64'h00ffffff00001000;

	lut_sub lut_2065 ({sk[592], i_2_, n_n95, n_n77, x108x, n_n953}, x153x);
	defparam lut_2065.LUT_SIZE = 6;
	defparam lut_2065.mask = 64'h00ffffff55575555;

	lut_sub lut_2068 ({sk[593], i_7_, i_8_, i_6_, x55x, n_n1052}, x263x);
	defparam lut_2068.LUT_SIZE = 6;
	defparam lut_2068.mask = 64'h00ffffff55555575;

	lut_sub lut_2071 ({sk[594], i_5_, i_3_, i_4_, n_n101, n_n83}, n_n975);
	defparam lut_2071.LUT_SIZE = 6;
	defparam lut_2071.mask = 64'h00ffffff00100000;

	lut_sub lut_2073 ({sk[595], i_7_, i_8_, i_6_, n_n84, n_n94}, n_n1184);
	defparam lut_2073.LUT_SIZE = 6;
	defparam lut_2073.mask = 64'h00ffffff00000001;

	lut_sub lut_2075 ({sk[596], i_7_, i_8_, i_6_, i_3_, i_4_}, x5493x);
	defparam lut_2075.LUT_SIZE = 6;
	defparam lut_2075.mask = 64'h00ffffff00001000;

	lut_sub lut_2077 ({sk[597], n_n93, n_n84, n_n102, n_n94, n_n85}, x224x);
	defparam lut_2077.LUT_SIZE = 6;
	defparam lut_2077.mask = 64'h00ffffff00000537;

	lut_sub lut_2080 ({sk[598], i_8_, i_6_, i_3_, x341x, n_n85}, x1384x);
	defparam lut_2080.LUT_SIZE = 6;
	defparam lut_2080.mask = 64'h00ffffff00000100;

	lut_sub lut_2082 ({sk[599], n_n91, n_n100, n_n102, x122x, x1008x}, x5599x);
	defparam lut_2082.LUT_SIZE = 6;
	defparam lut_2082.mask = 64'h00ffffff7777777f;

	lut_sub lut_2086 ({sk[600], n_n78, x252x, x43x, x49x, x348x}, x5600x);
	defparam lut_2086.LUT_SIZE = 6;
	defparam lut_2086.mask = 64'h00ffffff55ff7fff;

	lut_sub lut_2091 ({sk[601], n_n63, x41x, x234x, x242x, x5595x}, x5601x);
	defparam lut_2091.LUT_SIZE = 6;
	defparam lut_2091.mask = 64'h00ffffff575757ff;

	lut_sub lut_2095 ({sk[602], n_n1297, n_n1283, n_n1312, x309x, x326x}, x5602x);
	defparam lut_2095.LUT_SIZE = 6;
	defparam lut_2095.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2101 ({sk[603], n_n86, x104x, x21x, x123x, x217x}, x5603x);
	defparam lut_2101.LUT_SIZE = 6;
	defparam lut_2101.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_2106 ({sk[604], i_5_, i_3_, i_4_, n_n100}, x65x);
	defparam lut_2106.LUT_SIZE = 5;
	defparam lut_2106.mask = 32'h0f0f0001;

	lut_sub lut_2108 ({sk[605], i_5_, i_3_, i_4_, n_n82, n_n90}, x869x);
	defparam lut_2108.LUT_SIZE = 6;
	defparam lut_2108.mask = 64'h00ffffff00010000;

	lut_sub lut_2110 ({sk[606], n_n58, n_n95, x128x, x65x, x869x}, n_n211);
	defparam lut_2110.LUT_SIZE = 6;
	defparam lut_2110.mask = 64'h00ffffff55775f7f;

	lut_sub lut_2114 ({sk[607], x172x, n_n63, n_n85, x83x, x28x}, x120x);
	defparam lut_2114.LUT_SIZE = 6;
	defparam lut_2114.mask = 64'h00ffffff00330537;

	lut_sub lut_2117 ({sk[608], i_5_, i_3_, i_4_, n_n91, n_n83}, n_n1163);
	defparam lut_2117.LUT_SIZE = 6;
	defparam lut_2117.mask = 64'h00ffffff00100000;

	lut_sub lut_2119 ({sk[609], i_5_, i_3_, i_4_, n_n101, n_n83}, n_n1160);
	defparam lut_2119.LUT_SIZE = 6;
	defparam lut_2119.mask = 64'h00ffffff00000001;

	lut_sub lut_2121 ({sk[610], i_7_, i_8_, i_6_, n_n100, n_n84}, x1143x);
	defparam lut_2121.LUT_SIZE = 6;
	defparam lut_2121.mask = 64'h00ffffff00000010;

	lut_sub lut_2123 ({sk[611], i_5_, i_3_, i_4_, n_n101, n_n100}, n_n1216);
	defparam lut_2123.LUT_SIZE = 6;
	defparam lut_2123.mask = 64'h00ffffff01000000;

	lut_sub lut_2125 ({sk[612], i_7_, i_8_, i_6_, x63x}, n_n1158);
	defparam lut_2125.LUT_SIZE = 5;
	defparam lut_2125.mask = 32'h0f0f4000;

	lut_sub lut_2127 ({sk[613], i_5_, i_3_, i_4_, n_n101, n_n85}, n_n1146);
	defparam lut_2127.LUT_SIZE = 6;
	defparam lut_2127.mask = 64'h00ffffff00001000;

	lut_sub lut_2129 ({sk[614], i_7_, i_8_, i_6_, n_n84, n_n85}, n_n981);
	defparam lut_2129.LUT_SIZE = 6;
	defparam lut_2129.mask = 64'h00ffffff00000001;

	lut_sub lut_2131 ({sk[615], i_3_, i_4_, i_1_, i_0_, n_n93}, x617x);
	defparam lut_2131.LUT_SIZE = 6;
	defparam lut_2131.mask = 64'h00ffffff00001000;

	lut_sub lut_2133 ({sk[616], n_n74, n_n70, n_n63, n_n85, n_n40}, x5717x);
	defparam lut_2133.LUT_SIZE = 6;
	defparam lut_2133.mask = 64'h00ffffff00110313;

	lut_sub lut_2136 ({sk[617], i_3_, x341x, x37x, x139x, x6353x}, x5726x);
	defparam lut_2136.LUT_SIZE = 6;
	defparam lut_2136.mask = 64'h00ffffffbbbbbbbf;

	lut_sub lut_2140 ({sk[618], n_n91, x22x, n_n1181, x5715x, x6336x}, x5729x);
	defparam lut_2140.LUT_SIZE = 6;
	defparam lut_2140.mask = 64'h00ffffffbfbfbfff;

	lut_sub lut_2145 ({sk[619], n_n95, n_n1022, x237x, n_n1021, n_n994}, x5743x);
	defparam lut_2145.LUT_SIZE = 6;
	defparam lut_2145.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_2150 ({sk[620], i_3_, n_n1010, n_n1006, x313x, n_n1002}, x5744x);
	defparam lut_2150.LUT_SIZE = 6;
	defparam lut_2150.mask = 64'h00ffffff5fff7fff;

	lut_sub lut_2155 ({sk[621], n_n987, n_n984, x152x, x151x, x202x}, x5746x);
	defparam lut_2155.LUT_SIZE = 6;
	defparam lut_2155.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2161 ({sk[622], x188x, x114x, n_n296, x98x, x280x}, x6339x);
	defparam lut_2161.LUT_SIZE = 6;
	defparam lut_2161.mask = 64'h00ffffff80000000;

	lut_sub lut_2163 ({sk[623], i_5_, i_3_, i_4_, n_n101, n_n97}, n_n966);
	defparam lut_2163.LUT_SIZE = 6;
	defparam lut_2163.mask = 64'h00ffffff00010000;

	lut_sub lut_2165 ({sk[624], i_8_, i_6_, i_2_, n_n77, x175x}, x1017x);
	defparam lut_2165.LUT_SIZE = 6;
	defparam lut_2165.mask = 64'h00ffffff00000001;

	lut_sub lut_2167 ({sk[625], n_n91, n_n92, n_n100, n_n76, x129x}, x5392x);
	defparam lut_2167.LUT_SIZE = 6;
	defparam lut_2167.mask = 64'h00ffffff1111111f;

	lut_sub lut_2170 ({sk[626], i_2_, n_n101, n_n102, n_n942, x175x}, x79x);
	defparam lut_2170.LUT_SIZE = 6;
	defparam lut_2170.mask = 64'h00ffffff33333337;

	lut_sub lut_2173 ({sk[627], i_7_, i_8_, n_n40, n_n1057, n_n53}, x91x);
	defparam lut_2173.LUT_SIZE = 6;
	defparam lut_2173.mask = 64'h00ffffff33333337;

	lut_sub lut_2176 ({sk[628], i_3_, i_1_, i_2_, i_0_, x320x}, x103x);
	defparam lut_2176.LUT_SIZE = 6;
	defparam lut_2176.mask = 64'h00ffffff11000100;

	lut_sub lut_2179 ({sk[629], i_3_, n_n91, n_n85, x110x, n_n1108}, x161x);
	defparam lut_2179.LUT_SIZE = 6;
	defparam lut_2179.mask = 64'h00ffffff55555557;

	lut_sub lut_2182 ({sk[630], i_6_, x341x, n_n95, x34x, x85x}, x266x);
	defparam lut_2182.LUT_SIZE = 6;
	defparam lut_2182.mask = 64'h00ffffff03570303;

	lut_sub lut_2185 ({sk[631], i_7_, i_8_, i_6_, n_n1120, x128x}, x268x);
	defparam lut_2185.LUT_SIZE = 6;
	defparam lut_2185.mask = 64'h00ffffff33333733;

	lut_sub lut_2188 ({sk[632], i_5_, i_3_, i_4_, n_n78, n_n94}, n_n1177);
	defparam lut_2188.LUT_SIZE = 6;
	defparam lut_2188.mask = 64'h00ffffff00000010;

	lut_sub lut_2190 ({sk[633], i_7_, i_8_, n_n97, x127x, n_n1121}, x218x);
	defparam lut_2190.LUT_SIZE = 6;
	defparam lut_2190.mask = 64'h00ffffff55555755;

	lut_sub lut_2193 ({sk[634], n_n103, n_n82, n_n77, x107x, x218x}, x5826x);
	defparam lut_2193.LUT_SIZE = 6;
	defparam lut_2193.mask = 64'h00ffffff5757575f;

	lut_sub lut_2197 ({sk[635], i_6_, i_1_, i_0_, n_n58, x109x}, x526x);
	defparam lut_2197.LUT_SIZE = 6;
	defparam lut_2197.mask = 64'h00ffffff01000000;

	lut_sub lut_2199 ({sk[636], n_n63, n_n1153, x19x, x90x, x526x}, x5827x);
	defparam lut_2199.LUT_SIZE = 6;
	defparam lut_2199.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_2204 ({sk[637], n_n64, n_n52, x34x, n_n1047, x5835x}, x5841x);
	defparam lut_2204.LUT_SIZE = 6;
	defparam lut_2204.mask = 64'h00ffffff7777777f;

	lut_sub lut_2208 ({sk[638], n_n1105, x944x, x285x, x903x, x5492x}, x5842x);
	defparam lut_2208.LUT_SIZE = 6;
	defparam lut_2208.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2214 ({sk[639], n_n1109, n_n1095, x355x, n_n1088, x6335x}, x5844x);
	defparam lut_2214.LUT_SIZE = 6;
	defparam lut_2214.mask = 64'h00ffffffbfffffff;

	lut_sub lut_2220 ({sk[640], n_n1087, x805x, x263x, x161x, x102x}, x6334x);
	defparam lut_2220.LUT_SIZE = 6;
	defparam lut_2220.mask = 64'h00ffffff80000000;

	lut_sub lut_2222 ({sk[641], i_5_, i_3_, i_4_, i_2_, x108x}, x238x);
	defparam lut_2222.LUT_SIZE = 6;
	defparam lut_2222.mask = 64'h00ffffff04000000;

	lut_sub lut_2224 ({sk[642], i_7_, i_8_, i_6_, n_n1169, x238x}, x92x);
	defparam lut_2224.LUT_SIZE = 6;
	defparam lut_2224.mask = 64'h00ffffff33733333;

	lut_sub lut_2227 ({sk[643], n_n81, n_n101, n_n103, x38x, x322x}, x159x);
	defparam lut_2227.LUT_SIZE = 6;
	defparam lut_2227.mask = 64'h00ffffff1111111f;

	lut_sub lut_2230 ({sk[644], i_7_, i_8_, i_1_, i_2_, i_0_}, x247x);
	defparam lut_2230.LUT_SIZE = 6;
	defparam lut_2230.mask = 64'h00ffffff02000000;

	lut_sub lut_2232 ({sk[645], i_7_, i_8_, i_1_, i_2_, i_0_}, x316x);
	defparam lut_2232.LUT_SIZE = 6;
	defparam lut_2232.mask = 64'h00ffffff00000020;

	lut_sub lut_2234 ({sk[646], i_7_, i_8_, i_6_, n_n81, n_n97}, x335x);
	defparam lut_2234.LUT_SIZE = 6;
	defparam lut_2234.mask = 64'h00ffffff00001000;

	lut_sub lut_2236 ({sk[647], i_7_, i_8_, i_6_, n_n103, n_n84}, x344x);
	defparam lut_2236.LUT_SIZE = 6;
	defparam lut_2236.mask = 64'h00ffffff01000000;

	lut_sub lut_2238 ({sk[648], n_n73, x26x, n_n102, n_n1085, x20x}, x5886x);
	defparam lut_2238.LUT_SIZE = 6;
	defparam lut_2238.mask = 64'h00ffffff373737ff;

	lut_sub lut_2242 ({sk[649], n_n94, x334x, n_n1105, n_n1108, x5085x}, x5892x);
	defparam lut_2242.LUT_SIZE = 6;
	defparam lut_2242.mask = 64'h00ffffff3fff7fff;

	lut_sub lut_2247 ({sk[650], i_5_, i_3_, i_4_, n_n78, n_n100}, n_n1014);
	defparam lut_2247.LUT_SIZE = 6;
	defparam lut_2247.mask = 64'h00ffffff00000001;

	lut_sub lut_2249 ({sk[651], i_6_, n_n64, n_n85, x325x, x827x}, x152x);
	defparam lut_2249.LUT_SIZE = 6;
	defparam lut_2249.mask = 64'h00ffffff55555557;

	lut_sub lut_2252 ({sk[652], i_5_, i_3_, i_4_, n_n100, n_n95}, n_n1018);
	defparam lut_2252.LUT_SIZE = 6;
	defparam lut_2252.mask = 64'h00ffffff00000100;

	lut_sub lut_2254 ({sk[653], n_n91, x27x, n_n1074, n_n1045, n_n1060}, x5889x);
	defparam lut_2254.LUT_SIZE = 6;
	defparam lut_2254.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2259 ({sk[654], n_n1146, n_n1010, x5880x, x5881x, x5882x}, x5895x);
	defparam lut_2259.LUT_SIZE = 6;
	defparam lut_2259.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2265 ({sk[655], i_7_, i_8_, i_6_, x63x}, n_n999);
	defparam lut_2265.LUT_SIZE = 5;
	defparam lut_2265.mask = 32'h0f0f1000;

	lut_sub lut_2267 ({sk[656], i_7_, i_5_, i_6_, i_3_, n_n83}, x615x);
	defparam lut_2267.LUT_SIZE = 6;
	defparam lut_2267.mask = 64'h00ffffff00400000;

	lut_sub lut_2269 ({sk[657], n_n95, x44x, n_n980, n_n999, x615x}, x5901x);
	defparam lut_2269.LUT_SIZE = 6;
	defparam lut_2269.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2274 ({sk[658], n_n95, x29x, x829x, x125x, n_n947}, x5904x);
	defparam lut_2274.LUT_SIZE = 6;
	defparam lut_2274.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2279 ({sk[659], i_7_, i_8_, i_1_, i_2_, i_0_}, x129x);
	defparam lut_2279.LUT_SIZE = 6;
	defparam lut_2279.mask = 64'h00ffffff00040000;

	lut_sub lut_2281 ({sk[660], i_7_, i_8_, i_6_, x21x}, x877x);
	defparam lut_2281.LUT_SIZE = 5;
	defparam lut_2281.mask = 32'h0f0f0040;

	lut_sub lut_2283 ({sk[661], n_n93, x57x, x25x, n_n1177, x877x}, x5907x);
	defparam lut_2283.LUT_SIZE = 6;
	defparam lut_2283.mask = 64'h00ffffff77777fff;

	lut_sub lut_2288 ({sk[662], n_n52, n_n78, x34x, x52x, x22x}, x6361x);
	defparam lut_2288.LUT_SIZE = 6;
	defparam lut_2288.mask = 64'h00ffffff00770f7f;

	lut_sub lut_2296 ({sk[663], n_n78, n_n100, n_n84, n_n1216, x6361x}, x5908x);
	defparam lut_2296.LUT_SIZE = 6;
	defparam lut_2296.mask = 64'h00ffffff7777777f;

	lut_sub lut_2300 ({sk[664], n_n75, n_n81, n_n100, n_n40, x107x}, x155x);
	defparam lut_2300.LUT_SIZE = 6;
	defparam lut_2300.mask = 64'h00ffffff00550357;

	lut_sub lut_2303 ({sk[665], i_7_, i_8_, i_6_, n_n74, n_n90}, x332x);
	defparam lut_2303.LUT_SIZE = 6;
	defparam lut_2303.mask = 64'h00ffffff00000001;

	lut_sub lut_2305 ({sk[666], i_7_, i_8_, n_n54, n_n53, x332x}, x157x);
	defparam lut_2305.LUT_SIZE = 6;
	defparam lut_2305.mask = 64'h00ffffff55555755;

	lut_sub lut_2308 ({sk[667], i_3_, i_1_, i_2_}, x174x);
	defparam lut_2308.LUT_SIZE = 4;
	defparam lut_2308.mask = 16'h7704;

	lut_sub lut_2310 ({sk[668], i_7_, i_8_, n_n100, n_n1267, x131x}, x210x);
	defparam lut_2310.LUT_SIZE = 6;
	defparam lut_2310.mask = 64'h00ffffff33333337;

	lut_sub lut_2313 ({sk[669], i_5_, i_3_, i_4_, n_n78, n_n85}, x662x);
	defparam lut_2313.LUT_SIZE = 6;
	defparam lut_2313.mask = 64'h00ffffff00000010;

	lut_sub lut_2315 ({sk[670], i_1_, i_2_, i_0_, n_n101, n_n77}, x663x);
	defparam lut_2315.LUT_SIZE = 6;
	defparam lut_2315.mask = 64'h00ffffff00000010;

	lut_sub lut_2317 ({sk[671], i_7_, i_8_, i_6_, n_n84, n_n97}, x336x);
	defparam lut_2317.LUT_SIZE = 6;
	defparam lut_2317.mask = 64'h00ffffff00000001;

	lut_sub lut_2319 ({sk[672], i_5_, i_3_, i_4_, i_2_, x108x}, x33x);
	defparam lut_2319.LUT_SIZE = 6;
	defparam lut_2319.mask = 64'h00ffffff00100000;

	lut_sub lut_2321 ({sk[673], i_7_, i_8_, i_6_, x321x, x33x}, x226x);
	defparam lut_2321.LUT_SIZE = 6;
	defparam lut_2321.mask = 64'h00ffffff33333337;

	lut_sub lut_2324 ({sk[674], i_7_, i_8_, i_6_, n_n92, n_n100}, n_n1170);
	defparam lut_2324.LUT_SIZE = 6;
	defparam lut_2324.mask = 64'h00ffffff01000000;

	lut_sub lut_2326 ({sk[675], i_7_, i_8_, i_6_, x45x, x63x}, x267x);
	defparam lut_2326.LUT_SIZE = 6;
	defparam lut_2326.mask = 64'h00ffffff03050000;

	lut_sub lut_2329 ({sk[676], i_5_, i_6_, i_3_}, x130x);
	defparam lut_2329.LUT_SIZE = 4;
	defparam lut_2329.mask = 16'h7780;

	lut_sub lut_2331 ({sk[677], n_n93, n_n83, n_n102, x66x, x130x}, x5910x);
	defparam lut_2331.LUT_SIZE = 6;
	defparam lut_2331.mask = 64'h00ffffff1111111f;

	lut_sub lut_2334 ({sk[678], i_7_, i_8_, i_6_, x23x, x5910x}, x307x);
	defparam lut_2334.LUT_SIZE = 6;
	defparam lut_2334.mask = 64'h00ffffff55555575;

	lut_sub lut_2337 ({sk[679], i_7_, i_8_, i_3_}, x5686x);
	defparam lut_2337.LUT_SIZE = 4;
	defparam lut_2337.mask = 16'h7780;

	lut_sub lut_2339 ({sk[680], i_5_, i_6_, i_4_, i_1_, i_2_}, x5687x);
	defparam lut_2339.LUT_SIZE = 6;
	defparam lut_2339.mask = 64'h00ffffff00000200;

	lut_sub lut_2341 ({sk[681], i_7_, i_8_, i_6_, x42x}, n_n1164);
	defparam lut_2341.LUT_SIZE = 5;
	defparam lut_2341.mask = 32'h0f0f1000;

	lut_sub lut_2343 ({sk[682], i_5_, i_3_, i_4_, n_n91, n_n97}, n_n1088);
	defparam lut_2343.LUT_SIZE = 6;
	defparam lut_2343.mask = 64'h00ffffff00000010;

	lut_sub lut_2345 ({sk[683], i_5_, i_3_, i_4_, n_n101, n_n100}, x350x);
	defparam lut_2345.LUT_SIZE = 6;
	defparam lut_2345.mask = 64'h00ffffff00000100;

	lut_sub lut_2347 ({sk[684], i_7_, i_8_, n_n85, x348x, n_n40}, x5964x);
	defparam lut_2347.LUT_SIZE = 6;
	defparam lut_2347.mask = 64'h00ffffff33333733;

	lut_sub lut_2350 ({sk[685], n_n78, x323x, n_n1294, n_n1283, x22x}, x5975x);
	defparam lut_2350.LUT_SIZE = 6;
	defparam lut_2350.mask = 64'h00ffffff3fff7fff;

	lut_sub lut_2355 ({sk[686], x5965x, x5966x, x5967x, x5968x}, x5984x);
	defparam lut_2355.LUT_SIZE = 5;
	defparam lut_2355.mask = 32'h0f0f7fff;

	lut_sub lut_2360 ({sk[687], i_2_, n_n84, n_n70, n_n95, x108x}, x163x);
	defparam lut_2360.LUT_SIZE = 6;
	defparam lut_2360.mask = 64'h00ffffff00110005;

	lut_sub lut_2363 ({sk[688], i_5_, i_3_, i_4_, n_n83, n_n63}, n_n978);
	defparam lut_2363.LUT_SIZE = 6;
	defparam lut_2363.mask = 64'h00ffffff00000010;

	lut_sub lut_2365 ({sk[689], n_n91, n_n103, n_n102, x163x, n_n978}, x5990x);
	defparam lut_2365.LUT_SIZE = 6;
	defparam lut_2365.mask = 64'h00ffffff7777777f;

	lut_sub lut_2369 ({sk[690], n_n81, n_n101, n_n90, n_n999, x615x}, n_n296);
	defparam lut_2369.LUT_SIZE = 6;
	defparam lut_2369.mask = 64'h00ffffff7777777f;

	lut_sub lut_2373 ({sk[691], n_n100, n_n83, n_n74, n_n95, n_n296}, x5991x);
	defparam lut_2373.LUT_SIZE = 6;
	defparam lut_2373.mask = 64'h00ffffff55575757;

	lut_sub lut_2377 ({sk[692], i_3_, i_2_, i_0_}, x242x);
	defparam lut_2377.LUT_SIZE = 4;
	defparam lut_2377.mask = 16'h7702;

	lut_sub lut_2379 ({sk[693], i_1_, i_2_, i_0_, n_n91, n_n84}, x246x);
	defparam lut_2379.LUT_SIZE = 6;
	defparam lut_2379.mask = 64'h00ffffff00000010;

	lut_sub lut_2381 ({sk[694], i_5_, i_3_, i_4_, n_n101, n_n90}, x1557x);
	defparam lut_2381.LUT_SIZE = 6;
	defparam lut_2381.mask = 64'h00ffffff00000001;

	lut_sub lut_2383 ({sk[695], i_5_, i_3_, i_4_, n_n78, n_n97}, n_n1010);
	defparam lut_2383.LUT_SIZE = 6;
	defparam lut_2383.mask = 64'h00ffffff00100000;

	lut_sub lut_2385 ({sk[696], i_7_, i_8_, i_6_, x57x, x33x}, x270x);
	defparam lut_2385.LUT_SIZE = 6;
	defparam lut_2385.mask = 64'h00ffffff50300000;

	lut_sub lut_2388 ({sk[697], i_7_, i_5_, i_6_, n_n85, x54x}, n_n976);
	defparam lut_2388.LUT_SIZE = 6;
	defparam lut_2388.mask = 64'h00ffffff01000000;

	lut_sub lut_2390 ({sk[698], i_6_, i_3_, i_4_, x5068x, n_n976}, x272x);
	defparam lut_2390.LUT_SIZE = 6;
	defparam lut_2390.mask = 64'h00ffffff75555555;

	lut_sub lut_2393 ({sk[699], i_7_, i_8_, i_6_, x55x}, n_n1181);
	defparam lut_2393.LUT_SIZE = 5;
	defparam lut_2393.mask = 32'h0f0f4000;

	lut_sub lut_2395 ({sk[700], i_5_, i_3_, i_4_}, x194x);
	defparam lut_2395.LUT_SIZE = 4;
	defparam lut_2395.mask = 16'h7724;

	lut_sub lut_2398 ({sk[701], i_7_, i_8_, i_6_, n_n102, n_n97}, n_n987);
	defparam lut_2398.LUT_SIZE = 6;
	defparam lut_2398.mask = 64'h00ffffff01000000;

	lut_sub lut_2400 ({sk[702], i_7_, i_8_, i_6_, n_n103, n_n102}, n_n984);
	defparam lut_2400.LUT_SIZE = 6;
	defparam lut_2400.mask = 64'h00ffffff00100000;

	lut_sub lut_2402 ({sk[703], i_7_, i_8_, i_6_, x29x, x52x}, x147x);
	defparam lut_2402.LUT_SIZE = 6;
	defparam lut_2402.mask = 64'h00ffffff03500000;

	lut_sub lut_2405 ({sk[704], i_3_, x341x, n_n83, n_n82, n_n1021}, x274x);
	defparam lut_2405.LUT_SIZE = 6;
	defparam lut_2405.mask = 64'h00ffffff55555557;

	lut_sub lut_2408 ({sk[705], i_5_, i_3_, i_4_, n_n103, n_n95}, n_n1009);
	defparam lut_2408.LUT_SIZE = 6;
	defparam lut_2408.mask = 64'h00ffffff00000001;

	lut_sub lut_2410 ({sk[706], i_5_, i_6_, i_3_, n_n64, n_n103}, n_n1011);
	defparam lut_2410.LUT_SIZE = 6;
	defparam lut_2410.mask = 64'h00ffffff00000010;

	lut_sub lut_2412 ({sk[707], i_7_, i_8_, i_5_, i_6_, i_4_}, x339x);
	defparam lut_2412.LUT_SIZE = 6;
	defparam lut_2412.mask = 64'h00ffffff00800000;

	lut_sub lut_2414 ({sk[708], i_8_, i_6_, n_n81, x43x, x48x}, x217x);
	defparam lut_2414.LUT_SIZE = 6;
	defparam lut_2414.mask = 64'h00ffffff05053705;

	lut_sub lut_2417 ({sk[709], i_5_, n_n103, x54x, n_n82, x107x}, x71x);
	defparam lut_2417.LUT_SIZE = 6;
	defparam lut_2417.mask = 64'h00ffffff00000507;

	lut_sub lut_2420 ({sk[710], i_1_, i_2_, i_0_, n_n91, n_n102}, n_n994);
	defparam lut_2420.LUT_SIZE = 6;
	defparam lut_2420.mask = 64'h00ffffff00000010;

	lut_sub lut_2422 ({sk[711], i_1_, i_2_, i_0_, n_n74, n_n95}, n_n1006);
	defparam lut_2422.LUT_SIZE = 6;
	defparam lut_2422.mask = 64'h00ffffff00001000;

	lut_sub lut_2424 ({sk[712], i_7_, i_8_, n_n100, n_n54, n_n1006}, x59x);
	defparam lut_2424.LUT_SIZE = 6;
	defparam lut_2424.mask = 64'h00ffffff55555755;

	lut_sub lut_2427 ({sk[713], i_7_, i_6_, x109x, n_n982, n_n53}, x200x);
	defparam lut_2427.LUT_SIZE = 6;
	defparam lut_2427.mask = 64'h00ffffff33333733;

	lut_sub lut_2430 ({sk[714], i_1_, i_2_, i_0_, n_n38, n_n64}, x313x);
	defparam lut_2430.LUT_SIZE = 6;
	defparam lut_2430.mask = 64'h00ffffff00010000;

	lut_sub lut_2432 ({sk[715], i_8_, i_6_, n_n97, n_n947, x312x}, x5399x);
	defparam lut_2432.LUT_SIZE = 6;
	defparam lut_2432.mask = 64'h00ffffff33373333;

	lut_sub lut_2435 ({sk[716], i_7_, i_8_, i_6_, x76x}, n_n1013);
	defparam lut_2435.LUT_SIZE = 5;
	defparam lut_2435.mask = 32'h0f0f1000;

	lut_sub lut_2437 ({sk[717], i_1_, i_2_, i_0_, n_n63, n_n77}, n_n1028);
	defparam lut_2437.LUT_SIZE = 6;
	defparam lut_2437.mask = 64'h00ffffff00000001;

	lut_sub lut_2439 ({sk[718], i_5_, i_6_, i_4_, n_n86, n_n83}, x827x);
	defparam lut_2439.LUT_SIZE = 6;
	defparam lut_2439.mask = 64'h00ffffff00001000;

	lut_sub lut_2441 ({sk[719], i_7_, i_8_, i_2_, x108x, n_n76}, x753x);
	defparam lut_2441.LUT_SIZE = 6;
	defparam lut_2441.mask = 64'h00ffffff10000000;

	lut_sub lut_2443 ({sk[720], i_3_, i_2_, i_0_, x339x}, n_n1002);
	defparam lut_2443.LUT_SIZE = 5;
	defparam lut_2443.mask = 32'h0f0f0001;

	lut_sub lut_2445 ({sk[721], i_7_, i_8_, n_n74, n_n85, n_n1002}, x5609x);
	defparam lut_2445.LUT_SIZE = 6;
	defparam lut_2445.mask = 64'h00ffffff55555557;

	lut_sub lut_2448 ({sk[722], i_6_, n_n86, x112x, n_n1001, x152x}, x5616x);
	defparam lut_2448.LUT_SIZE = 6;
	defparam lut_2448.mask = 64'h00ffffff7777777f;

	lut_sub lut_2452 ({sk[723], x25x, n_n82, n_n1047, n_n1013, n_n1014}, x5617x);
	defparam lut_2452.LUT_SIZE = 6;
	defparam lut_2452.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2457 ({sk[724], n_n980, n_n983, n_n986, n_n1021, n_n1028}, x5618x);
	defparam lut_2457.LUT_SIZE = 6;
	defparam lut_2457.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2463 ({sk[725], n_n86, n_n85, n_n76, x5609x, x299x}, x5619x);
	defparam lut_2463.LUT_SIZE = 6;
	defparam lut_2463.mask = 64'h00ffffff7777777f;

	lut_sub lut_2467 ({sk[726], n_n78, x29x, x201x, x271x, x275x}, x5620x);
	defparam lut_2467.LUT_SIZE = 6;
	defparam lut_2467.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2472 ({sk[727], i_7_, i_8_, i_6_, x21x}, x345x);
	defparam lut_2472.LUT_SIZE = 5;
	defparam lut_2472.mask = 32'h0f0f0001;

	lut_sub lut_2474 ({sk[728], i_7_, i_6_, i_3_, x341x, n_n97}, x249x);
	defparam lut_2474.LUT_SIZE = 6;
	defparam lut_2474.mask = 64'h00ffffff00000001;

	lut_sub lut_2476 ({sk[729], i_7_, i_8_, i_5_, i_6_, n_n83}, x1583x);
	defparam lut_2476.LUT_SIZE = 6;
	defparam lut_2476.mask = 64'h00ffffff10000000;

	lut_sub lut_2478 ({sk[730], i_3_, i_1_, i_0_, n_n70, n_n71}, n_n1026);
	defparam lut_2478.LUT_SIZE = 6;
	defparam lut_2478.mask = 64'h00ffffff00100000;

	lut_sub lut_2480 ({sk[731], i_7_, i_8_, i_6_, i_4_}, x4876x);
	defparam lut_2480.LUT_SIZE = 5;
	defparam lut_2480.mask = 32'h0f0f0080;

	lut_sub lut_2482 ({sk[732], i_7_, i_6_, i_3_, i_4_, n_n85}, x1581x);
	defparam lut_2482.LUT_SIZE = 6;
	defparam lut_2482.mask = 64'h00ffffff00001000;

	lut_sub lut_2484 ({sk[733], i_1_, x56x, n_n1026, x4876x, x1581x}, x288x);
	defparam lut_2484.LUT_SIZE = 6;
	defparam lut_2484.mask = 64'h00ffffff5f5f5f7f;

	lut_sub lut_2488 ({sk[734], i_7_, i_8_, i_6_, n_n92, n_n90}, n_n943);
	defparam lut_2488.LUT_SIZE = 6;
	defparam lut_2488.mask = 64'h00ffffff01000000;

	lut_sub lut_2490 ({sk[735], i_2_, n_n81, n_n91, n_n82, x175x}, x202x);
	defparam lut_2490.LUT_SIZE = 6;
	defparam lut_2490.mask = 64'h00ffffff00050011;

	lut_sub lut_2493 ({sk[736], i_7_, i_2_, x108x, n_n76, n_n1004}, x203x);
	defparam lut_2493.LUT_SIZE = 6;
	defparam lut_2493.mask = 64'h00ffffff55575555;

	lut_sub lut_2496 ({sk[737], i_0_, n_n91, x75x, n_n77, x34x}, x225x);
	defparam lut_2496.LUT_SIZE = 6;
	defparam lut_2496.mask = 64'h00ffffff00550057;

	lut_sub lut_2499 ({sk[738], i_5_, i_3_, i_4_, n_n93, n_n85}, x1008x);
	defparam lut_2499.LUT_SIZE = 6;
	defparam lut_2499.mask = 64'h00ffffff10000000;

	lut_sub lut_2501 ({sk[739], n_n81, n_n91, x41x, x20x, x1008x}, x289x);
	defparam lut_2501.LUT_SIZE = 6;
	defparam lut_2501.mask = 64'h00ffffff555f777f;

	lut_sub lut_2505 ({sk[740], i_5_, i_3_, i_4_, n_n78, n_n90}, x1153x);
	defparam lut_2505.LUT_SIZE = 6;
	defparam lut_2505.mask = 64'h00ffffff00010000;

	lut_sub lut_2507 ({sk[741], n_n93, n_n102, n_n63, n_n77, n_n90}, x5407x);
	defparam lut_2507.LUT_SIZE = 6;
	defparam lut_2507.mask = 64'h00ffffff00051115;

	lut_sub lut_2510 ({sk[742], i_3_, n_n52, n_n83, x109x, n_n1009}, x98x);
	defparam lut_2510.LUT_SIZE = 6;
	defparam lut_2510.mask = 64'h00ffffff55575555;

	lut_sub lut_2513 ({sk[743], i_3_, i_4_, n_n38, n_n103, n_n1043}, x154x);
	defparam lut_2513.LUT_SIZE = 6;
	defparam lut_2513.mask = 64'h00ffffff57555555;

	lut_sub lut_2516 ({sk[744], i_3_, i_0_, n_n101, x75x, n_n1022}, x212x);
	defparam lut_2516.LUT_SIZE = 6;
	defparam lut_2516.mask = 64'h00ffffff55575555;

	lut_sub lut_2519 ({sk[745], i_8_, i_6_, n_n102, n_n94, n_n1028}, x280x);
	defparam lut_2519.LUT_SIZE = 6;
	defparam lut_2519.mask = 64'h00ffffff55575555;

	lut_sub lut_2522 ({sk[746], n_n94, n_n1010, x5085x, x249x, n_n1026}, x5791x);
	defparam lut_2522.LUT_SIZE = 6;
	defparam lut_2522.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_2527 ({sk[747], n_n1032, n_n1040, x114x, n_n1011, x59x}, x5792x);
	defparam lut_2527.LUT_SIZE = 6;
	defparam lut_2527.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2533 ({sk[748], n_n1046, x274x, x151x, x1583x, x98x}, x5793x);
	defparam lut_2533.LUT_SIZE = 6;
	defparam lut_2533.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2539 ({sk[749], n_n1045, n_n1013, x154x, x212x, x280x}, x6333x);
	defparam lut_2539.LUT_SIZE = 6;
	defparam lut_2539.mask = 64'h00ffffff80000000;

	lut_sub lut_2541 ({sk[750], i_7_, i_8_, i_6_, x58x, x44x}, x101x);
	defparam lut_2541.LUT_SIZE = 6;
	defparam lut_2541.mask = 64'h00ffffff00503000;

	lut_sub lut_2544 ({sk[751], i_5_, i_3_, n_n93, n_n97, x900x}, x102x);
	defparam lut_2544.LUT_SIZE = 6;
	defparam lut_2544.mask = 64'h00ffffff55555557;

	lut_sub lut_2547 ({sk[752], n_n91, n_n84, n_n85, n_n1108, x92x}, x5504x);
	defparam lut_2547.LUT_SIZE = 6;
	defparam lut_2547.mask = 64'h00ffffff7777777f;

	lut_sub lut_2551 ({sk[753], n_n86, n_n97, n_n77, n_n1128, x224x}, x5505x);
	defparam lut_2551.LUT_SIZE = 6;
	defparam lut_2551.mask = 64'h00ffffff7777777f;

	lut_sub lut_2555 ({sk[754], n_n38, n_n64, x64x, n_n1132, x5499x}, x5507x);
	defparam lut_2555.LUT_SIZE = 6;
	defparam lut_2555.mask = 64'h00ffffff7777777f;

	lut_sub lut_2559 ({sk[755], i_7_, i_8_, i_6_, n_n81, n_n103}, x876x);
	defparam lut_2559.LUT_SIZE = 6;
	defparam lut_2559.mask = 64'h00ffffff01000000;

	lut_sub lut_2561 ({sk[756], i_0_, x75x, n_n82, n_n95, n_n77}, x166x);
	defparam lut_2561.LUT_SIZE = 6;
	defparam lut_2561.mask = 64'h00ffffff00110005;

	lut_sub lut_2564 ({sk[757], i_7_, i_8_, n_n74, x20x, x65x}, x220x);
	defparam lut_2564.LUT_SIZE = 6;
	defparam lut_2564.mask = 64'h00ffffff03035703;

	lut_sub lut_2567 ({sk[758], i_3_, x341x, n_n78, n_n97, n_n1172}, x281x);
	defparam lut_2567.LUT_SIZE = 6;
	defparam lut_2567.mask = 64'h00ffffff55555557;

	lut_sub lut_2570 ({sk[759], i_7_, i_8_, i_6_, x45x, x239x}, x5514x);
	defparam lut_2570.LUT_SIZE = 6;
	defparam lut_2570.mask = 64'h00ffffff00050300;

	lut_sub lut_2573 ({sk[760], n_n74, x662x, x663x, x31x, x1153x}, x5699x);
	defparam lut_2573.LUT_SIZE = 6;
	defparam lut_2573.mask = 64'h00ffffff5fff7fff;

	lut_sub lut_2578 ({sk[761], n_n91, x42x, n_n1259, x344x, n_n1312}, x5700x);
	defparam lut_2578.LUT_SIZE = 6;
	defparam lut_2578.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2583 ({sk[762], n_n101, n_n91, x33x, x65x, x5697x}, x5703x);
	defparam lut_2583.LUT_SIZE = 6;
	defparam lut_2583.mask = 64'h00ffffff55775f7f;

	lut_sub lut_2587 ({sk[763], x104x, x157x, x289x}, x5704x);
	defparam lut_2587.LUT_SIZE = 4;
	defparam lut_2587.mask = 16'h777f;

	lut_sub lut_2591 ({sk[764], x343x, n_n1215, x5693x, x5694x, x5695x}, x5706x);
	defparam lut_2591.LUT_SIZE = 6;
	defparam lut_2591.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2597 ({sk[765], i_7_, i_8_, i_0_, x75x, n_n66}, x1508x);
	defparam lut_2597.LUT_SIZE = 6;
	defparam lut_2597.mask = 64'h00ffffff00010000;

	lut_sub lut_2599 ({sk[766], i_5_, i_3_, n_n93, n_n85, x1508x}, x121x);
	defparam lut_2599.LUT_SIZE = 6;
	defparam lut_2599.mask = 64'h00ffffff55555755;

	lut_sub lut_2602 ({sk[767], i_8_, i_6_, n_n92, n_n97, x68x}, x287x);
	defparam lut_2602.LUT_SIZE = 6;
	defparam lut_2602.mask = 64'h00ffffff55575555;

	lut_sub lut_2605 ({sk[768], i_3_, x45x, x110x, x331x, x316x}, x122x);
	defparam lut_2605.LUT_SIZE = 6;
	defparam lut_2605.mask = 64'h00ffffff05370033;

	lut_sub lut_2608 ({sk[769], i_7_, i_8_, i_2_, x175x, n_n66}, x900x);
	defparam lut_2608.LUT_SIZE = 6;
	defparam lut_2608.mask = 64'h00ffffff00000010;

	lut_sub lut_2610 ({sk[770], i_5_, i_3_, i_4_, n_n93, n_n94}, x1440x);
	defparam lut_2610.LUT_SIZE = 6;
	defparam lut_2610.mask = 64'h00ffffff00100000;

	lut_sub lut_2612 ({sk[771], i_3_, i_4_}, x312x);
	defparam lut_2612.LUT_SIZE = 3;
	defparam lut_2612.mask = 8'h52;

	lut_sub lut_2614 ({sk[772], i_7_, i_8_, i_0_}, x5828x);
	defparam lut_2614.LUT_SIZE = 4;
	defparam lut_2614.mask = 16'h7704;

	lut_sub lut_2616 ({sk[773], i_7_, i_8_, i_6_, x57x}, x670x);
	defparam lut_2616.LUT_SIZE = 5;
	defparam lut_2616.mask = 32'h0f0f0010;

	lut_sub lut_2618 ({sk[774], i_5_, i_3_, i_4_, n_n94, n_n95}, x835x);
	defparam lut_2618.LUT_SIZE = 6;
	defparam lut_2618.mask = 64'h00ffffff00000001;

	lut_sub lut_2620 ({sk[775], i_7_, i_6_, i_3_, n_n83, x109x}, x1085x);
	defparam lut_2620.LUT_SIZE = 6;
	defparam lut_2620.mask = 64'h00ffffff00000010;

	lut_sub lut_2622 ({sk[776], i_5_, i_6_, i_3_, n_n64, n_n90}, x1108x);
	defparam lut_2622.LUT_SIZE = 6;
	defparam lut_2622.mask = 64'h00ffffff00000001;

	lut_sub lut_2624 ({sk[777], i_8_, i_5_, i_1_, n_n52, x56x}, x1442x);
	defparam lut_2624.LUT_SIZE = 6;
	defparam lut_2624.mask = 64'h00ffffff00000001;

	lut_sub lut_2626 ({sk[778], i_7_, i_8_, i_5_, i_6_, n_n100}, x1446x);
	defparam lut_2626.LUT_SIZE = 6;
	defparam lut_2626.mask = 64'h00ffffff04000000;

	lut_sub lut_2628 ({sk[779], i_7_, i_8_, i_6_, n_n81, x75x}, x1589x);
	defparam lut_2628.LUT_SIZE = 6;
	defparam lut_2628.mask = 64'h00ffffff00010000;

	lut_sub lut_2630 ({sk[780], n_n81, n_n52, x172x, n_n85, x311x}, x4848x);
	defparam lut_2630.LUT_SIZE = 6;
	defparam lut_2630.mask = 64'h00ffffff05050537;

	lut_sub lut_2633 ({sk[781], i_7_, i_8_, i_6_, x27x, x45x}, x4849x);
	defparam lut_2633.LUT_SIZE = 6;
	defparam lut_2633.mask = 64'h00ffffff00700700;

	lut_sub lut_2638 ({sk[782], n_n101, n_n78, n_n74, n_n97, x55x}, x4852x);
	defparam lut_2638.LUT_SIZE = 6;
	defparam lut_2638.mask = 64'h00ffffff00035557;

	lut_sub lut_2641 ({sk[783], n_n93, x57x, x26x, x235x, x329x}, x4858x);
	defparam lut_2641.LUT_SIZE = 6;
	defparam lut_2641.mask = 64'h00ffffff77777fff;

	lut_sub lut_2646 ({sk[784], n_n52, n_n93, x64x, x112x, x4849x}, x4860x);
	defparam lut_2646.LUT_SIZE = 6;
	defparam lut_2646.mask = 64'h00ffffff555f777f;

	lut_sub lut_2650 ({sk[785], n_n81, n_n64, n_n52, n_n103, n_n1011}, x4885x);
	defparam lut_2650.LUT_SIZE = 6;
	defparam lut_2650.mask = 64'h00ffffff55555557;

	lut_sub lut_2653 ({sk[786], x55x, n_n95, n_n1043, n_n1059, n_n1042}, x6348x);
	defparam lut_2653.LUT_SIZE = 6;
	defparam lut_2653.mask = 64'h00ffffff80808000;

	lut_sub lut_2656 ({sk[787], n_n75, n_n81, n_n93, n_n103, n_n77}, x4935x);
	defparam lut_2656.LUT_SIZE = 6;
	defparam lut_2656.mask = 64'h00ffffff01010133;

	lut_sub lut_2659 ({sk[788], n_n81, n_n86, n_n91, x64x, x108x}, x4961x);
	defparam lut_2659.LUT_SIZE = 6;
	defparam lut_2659.mask = 64'h00ffffff03030357;

	lut_sub lut_2662 ({sk[789], i_1_, i_2_, n_n58, n_n102, x1446x}, x4967x);
	defparam lut_2662.LUT_SIZE = 6;
	defparam lut_2662.mask = 64'h00ffffff55555557;

	lut_sub lut_2665 ({sk[790], i_5_, i_6_, x54x, x37x, x328x}, x4968x);
	defparam lut_2665.LUT_SIZE = 6;
	defparam lut_2665.mask = 64'h00ffffff03070005;

	lut_sub lut_2668 ({sk[791], i_3_, x27x, n_n97, n_n82, x325x}, x4969x);
	defparam lut_2668.LUT_SIZE = 6;
	defparam lut_2668.mask = 64'h00ffffff00330133;

	lut_sub lut_2671 ({sk[792], n_n73, n_n92, n_n103, n_n82, n_n77}, x4970x);
	defparam lut_2671.LUT_SIZE = 6;
	defparam lut_2671.mask = 64'h00ffffff0101010f;

	lut_sub lut_2674 ({sk[793], n_n80, n_n86, x105x, x109x, x1442x}, x4971x);
	defparam lut_2674.LUT_SIZE = 6;
	defparam lut_2674.mask = 64'h00ffffff5f5f5f7f;

	lut_sub lut_2678 ({sk[794], i_7_, i_6_, n_n1082, x207x, x21x}, x4972x);
	defparam lut_2678.LUT_SIZE = 6;
	defparam lut_2678.mask = 64'h00ffffff7f3f3f3f;

	lut_sub lut_2682 ({sk[795], i_7_, i_8_, x254x, x53x, x63x}, x4973x);
	defparam lut_2682.LUT_SIZE = 6;
	defparam lut_2682.mask = 64'h00ffffff0f5f3f0f;

	lut_sub lut_2686 ({sk[796], n_n81, n_n95, n_n1078, n_n90, x4961x}, x4974x);
	defparam lut_2686.LUT_SIZE = 6;
	defparam lut_2686.mask = 64'h00ffffff5f5f5f7f;

	lut_sub lut_2690 ({sk[797], x245x, x38x, n_n1279, n_n1153, n_n1297}, x4975x);
	defparam lut_2690.LUT_SIZE = 6;
	defparam lut_2690.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2695 ({sk[798], n_n91, x27x, n_n1324, x251x, x321x}, x4976x);
	defparam lut_2695.LUT_SIZE = 6;
	defparam lut_2695.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2700 ({sk[799], x4967x, x4968x, x4969x, x4970x}, x4982x);
	defparam lut_2700.LUT_SIZE = 5;
	defparam lut_2700.mask = 32'h0f0f7fff;

	lut_sub lut_2705 ({sk[800], i_7_, i_8_, i_6_, x21x, x34x}, x5035x);
	defparam lut_2705.LUT_SIZE = 6;
	defparam lut_2705.mask = 64'h00ffffff33500000;

	lut_sub lut_2708 ({sk[801], n_n93, n_n74, n_n97, n_n1188, x178x}, x5037x);
	defparam lut_2708.LUT_SIZE = 6;
	defparam lut_2708.mask = 64'h00ffffff7777777f;

	lut_sub lut_2712 ({sk[802], n_n38, n_n70, x34x, x354x, x62x}, x5056x);
	defparam lut_2712.LUT_SIZE = 6;
	defparam lut_2712.mask = 64'h00ffffff1111111f;

	lut_sub lut_2715 ({sk[803], n_n93, n_n1185, n_n1172, x19x, x36x}, x5059x);
	defparam lut_2715.LUT_SIZE = 6;
	defparam lut_2715.mask = 64'h00ffffff0fff7fff;

	lut_sub lut_2720 ({sk[804], i_7_, i_8_, i_6_, x64x, x53x}, x5087x);
	defparam lut_2720.LUT_SIZE = 6;
	defparam lut_2720.mask = 64'h00ffffff00000070;

	lut_sub lut_2723 ({sk[805], n_n52, n_n101, x39x, x58x, x1359x}, x5093x);
	defparam lut_2723.LUT_SIZE = 6;
	defparam lut_2723.mask = 64'h00ffffff55775f7f;

	lut_sub lut_2727 ({sk[806], x337x, n_n1039, n_n1091, x322x, n_n1103}, x5099x);
	defparam lut_2727.LUT_SIZE = 6;
	defparam lut_2727.mask = 64'h00ffffff5fff7fff;

	lut_sub lut_2732 ({sk[807], x49x, n_n1120, n_n1052, n_n1331, x177x}, x5100x);
	defparam lut_2732.LUT_SIZE = 6;
	defparam lut_2732.mask = 64'h00ffffff3fff7fff;

	lut_sub lut_2737 ({sk[808], n_n82, x21x, x46x, x173x, x233x}, x5101x);
	defparam lut_2737.LUT_SIZE = 6;
	defparam lut_2737.mask = 64'h00ffffff55775f7f;

	lut_sub lut_2741 ({sk[809], x117x, x133x, x148x, x323x, x1352x}, x5103x);
	defparam lut_2741.LUT_SIZE = 6;
	defparam lut_2741.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2747 ({sk[810], n_n83, x35x, x201x, x256x, x271x}, x5104x);
	defparam lut_2747.LUT_SIZE = 6;
	defparam lut_2747.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2752 ({sk[811], i_3_, x341x, n_n83, n_n82, n_n989}, x5114x);
	defparam lut_2752.LUT_SIZE = 6;
	defparam lut_2752.mask = 64'h00ffffff55555557;

	lut_sub lut_2755 ({sk[812], n_n64, n_n101, n_n85, x49x, n_n76}, x5148x);
	defparam lut_2755.LUT_SIZE = 6;
	defparam lut_2755.mask = 64'h00ffffff00330537;

	lut_sub lut_2758 ({sk[813], x27x, x113x, n_n63, n_n95, x34x}, x5150x);
	defparam lut_2758.LUT_SIZE = 6;
	defparam lut_2758.mask = 64'h00ffffff05ff37ff;

	lut_sub lut_2762 ({sk[814], n_n101, n_n83, n_n102, x105x, x1359x}, x5151x);
	defparam lut_2762.LUT_SIZE = 6;
	defparam lut_2762.mask = 64'h00ffffff7777777f;

	lut_sub lut_2766 ({sk[815], n_n101, n_n103, n_n84, x117x, x1292x}, x5152x);
	defparam lut_2766.LUT_SIZE = 6;
	defparam lut_2766.mask = 64'h00ffffff7777777f;

	lut_sub lut_2770 ({sk[816], n_n93, n_n84, x233x, x36x, x48x}, x5159x);
	defparam lut_2770.LUT_SIZE = 6;
	defparam lut_2770.mask = 64'h00ffffff0f5f3f7f;

	lut_sub lut_2774 ({sk[817], i_7_, i_8_, i_6_, x352x, x63x}, x5205x);
	defparam lut_2774.LUT_SIZE = 6;
	defparam lut_2774.mask = 64'h00ffffff33333733;

	lut_sub lut_2777 ({sk[818], i_2_, n_n91, x56x, x49x, x318x}, x5206x);
	defparam lut_2777.LUT_SIZE = 6;
	defparam lut_2777.mask = 64'h00ffffff05370033;

	lut_sub lut_2780 ({sk[819], i_7_, i_8_, i_6_, x105x, x41x}, x5208x);
	defparam lut_2780.LUT_SIZE = 6;
	defparam lut_2780.mask = 64'h00ffffff37333333;

	lut_sub lut_2783 ({sk[820], i_7_, i_8_, i_6_, x46x, x5206x}, x5214x);
	defparam lut_2783.LUT_SIZE = 6;
	defparam lut_2783.mask = 64'h00ffffff55557557;

	lut_sub lut_2787 ({sk[821], x323x, n_n1330, x185x, x258x, x5205x}, x5217x);
	defparam lut_2787.LUT_SIZE = 6;
	defparam lut_2787.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2793 ({sk[822], n_n77, x1291x, x1292x, x183x, x31x}, x6355x);
	defparam lut_2793.LUT_SIZE = 6;
	defparam lut_2793.mask = 64'h00ffffffc0008000;

	lut_sub lut_2796 ({sk[823], n_n78, x67x, n_n1057, n_n1125, x248x}, x5244x);
	defparam lut_2796.LUT_SIZE = 6;
	defparam lut_2796.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2801 ({sk[824], i_8_, x341x, n_n52, x75x, x252x}, x5283x);
	defparam lut_2801.LUT_SIZE = 6;
	defparam lut_2801.mask = 64'h00ffffff55555557;

	lut_sub lut_2804 ({sk[825], i_1_, n_n64, n_n40, x30x, x1108x}, x5288x);
	defparam lut_2804.LUT_SIZE = 6;
	defparam lut_2804.mask = 64'h00ffffff55555557;

	lut_sub lut_2807 ({sk[826], i_1_, i_2_, n_n70, n_n77, n_n87}, x6356x);
	defparam lut_2807.LUT_SIZE = 6;
	defparam lut_2807.mask = 64'h00fffffffffeffff;

	lut_sub lut_2819 ({sk[827], i_7_, i_8_, i_4_, x311x, x6356x}, x5289x);
	defparam lut_2819.LUT_SIZE = 6;
	defparam lut_2819.mask = 64'h00ffffffaaabaaaa;

	lut_sub lut_2822 ({sk[828], n_n93, n_n102, x127x, x328x, x175x}, x5290x);
	defparam lut_2822.LUT_SIZE = 6;
	defparam lut_2822.mask = 64'h00ffffff03030357;

	lut_sub lut_2825 ({sk[829], i_7_, i_8_, n_n103, n_n100, n_n76}, x5291x);
	defparam lut_2825.LUT_SIZE = 6;
	defparam lut_2825.mask = 64'h00ffffff05000011;

	lut_sub lut_2828 ({sk[830], i_4_, x234x, x66x, x242x, x28x}, x5292x);
	defparam lut_2828.LUT_SIZE = 6;
	defparam lut_2828.mask = 64'h00ffffff05370033;

	lut_sub lut_2831 ({sk[831], n_n93, n_n84, x109x, n_n90, x85x}, x5293x);
	defparam lut_2831.LUT_SIZE = 6;
	defparam lut_2831.mask = 64'h00ffffff05050537;

	lut_sub lut_2834 ({sk[832], n_n91, x58x, n_n82, x67x, x5293x}, x5305x);
	defparam lut_2834.LUT_SIZE = 6;
	defparam lut_2834.mask = 64'h00ffffff555f777f;

	lut_sub lut_2838 ({sk[833], i_7_, i_8_, x32x, n_n74, x44x}, x6349x);
	defparam lut_2838.LUT_SIZE = 6;
	defparam lut_2838.mask = 64'h00ffffffa8fcfcfc;

	lut_sub lut_2845 ({sk[834], n_n1217, x174x, x336x, x246x, x339x}, x6346x);
	defparam lut_2845.LUT_SIZE = 6;
	defparam lut_2845.mask = 64'h00ffffffc0800000;

	lut_sub lut_2848 ({sk[835], i_8_, i_6_, i_3_, n_n85, n_n1030}, x5321x);
	defparam lut_2848.LUT_SIZE = 6;
	defparam lut_2848.mask = 64'h00ffffff75555555;

	lut_sub lut_2851 ({sk[836], i_7_, i_8_, i_6_, x55x, n_n1058}, x5322x);
	defparam lut_2851.LUT_SIZE = 6;
	defparam lut_2851.mask = 64'h00ffffff55555557;

	lut_sub lut_2854 ({sk[837], i_1_, i_2_, n_n64, x109x, x83x}, x5342x);
	defparam lut_2854.LUT_SIZE = 6;
	defparam lut_2854.mask = 64'h00ffffff55555557;

	lut_sub lut_2857 ({sk[838], i_6_, n_n70, x110x, n_n53, x319x}, x5351x);
	defparam lut_2857.LUT_SIZE = 6;
	defparam lut_2857.mask = 64'h00ffffff55575555;

	lut_sub lut_2860 ({sk[839], n_n101, n_n989, x52x, n_n944, n_n982}, x5358x);
	defparam lut_2860.LUT_SIZE = 6;
	defparam lut_2860.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_2865 ({sk[840], n_n78, x42x, n_n967, n_n1121, x236x}, x5359x);
	defparam lut_2865.LUT_SIZE = 6;
	defparam lut_2865.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2870 ({sk[841], n_n73, x42x, x111x, x5342x, x5351x}, x5360x);
	defparam lut_2870.LUT_SIZE = 6;
	defparam lut_2870.mask = 64'h00ffffff7777777f;

	lut_sub lut_2874 ({sk[842], n_n101, x97x, x145x, n_n951, x44x}, x5362x);
	defparam lut_2874.LUT_SIZE = 6;
	defparam lut_2874.mask = 64'h00ffffff3fff7fff;

	lut_sub lut_2879 ({sk[843], i_8_, x70x, x215x, x262x, x275x}, x5364x);
	defparam lut_2879.LUT_SIZE = 6;
	defparam lut_2879.mask = 64'h00ffffff7fff7f7f;

	lut_sub lut_2884 ({sk[844], x245x, x38x, n_n1093, n_n1074, n_n1087}, x6344x);
	defparam lut_2884.LUT_SIZE = 6;
	defparam lut_2884.mask = 64'h00ffffff80808000;

	lut_sub lut_2887 ({sk[845], n_n80, n_n83, x234x, x320x, n_n973}, x6351x);
	defparam lut_2887.LUT_SIZE = 6;
	defparam lut_2887.mask = 64'h00ffffffaa88a080;

	lut_sub lut_2892 ({sk[846], i_3_, n_n78, n_n85, x37x, x109x}, x5411x);
	defparam lut_2892.LUT_SIZE = 6;
	defparam lut_2892.mask = 64'h00ffffff00001115;

	lut_sub lut_2895 ({sk[847], n_n70, x48x, n_n87, x194x, x353x}, x5429x);
	defparam lut_2895.LUT_SIZE = 6;
	defparam lut_2895.mask = 64'h00ffffff00330537;

	lut_sub lut_2898 ({sk[848], i_5_, i_6_, n_n75, x251x, n_n90}, x5446x);
	defparam lut_2898.LUT_SIZE = 6;
	defparam lut_2898.mask = 64'h00ffffff33373333;

	lut_sub lut_2901 ({sk[849], i_7_, i_3_, n_n1078, n_n40, x330x}, x5460x);
	defparam lut_2901.LUT_SIZE = 6;
	defparam lut_2901.mask = 64'h00ffffff0f0f0f1f;

	lut_sub lut_2904 ({sk[850], i_8_, i_2_, n_n54, x56x, x355x}, x5467x);
	defparam lut_2904.LUT_SIZE = 6;
	defparam lut_2904.mask = 64'h00ffffff55555755;

	lut_sub lut_2907 ({sk[851], i_8_, n_n85, x127x, x21x, x173x}, x5468x);
	defparam lut_2907.LUT_SIZE = 6;
	defparam lut_2907.mask = 64'h00ffffff1111111f;

	lut_sub lut_2910 ({sk[852], i_7_, i_6_, x26x, n_n1085, x279x}, x5472x);
	defparam lut_2910.LUT_SIZE = 6;
	defparam lut_2910.mask = 64'h00ffffff7f777777;

	lut_sub lut_2914 ({sk[853], i_6_, n_n86, x43x, n_n1125, x5460x}, x5474x);
	defparam lut_2914.LUT_SIZE = 6;
	defparam lut_2914.mask = 64'h00ffffff7777777f;

	lut_sub lut_2918 ({sk[854], n_n73, n_n1082, x36x, n_n1045, n_n1043}, x5475x);
	defparam lut_2918.LUT_SIZE = 6;
	defparam lut_2918.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_2923 ({sk[855], n_n91, n_n40, x66x, x44x, x5468x}, x5478x);
	defparam lut_2923.LUT_SIZE = 6;
	defparam lut_2923.mask = 64'h00ffffff555f777f;

	lut_sub lut_2927 ({sk[856], x141x, x142x, x150x, n_n1046, n_n1047}, x5479x);
	defparam lut_2927.LUT_SIZE = 6;
	defparam lut_2927.mask = 64'h00ffffff7fffffff;

	lut_sub lut_2933 ({sk[857], n_n1118, n_n1030, x66x, x5442x, n_n1101}, x6343x);
	defparam lut_2933.LUT_SIZE = 6;
	defparam lut_2933.mask = 64'h00ffffffa8000000;

	lut_sub lut_2936 ({sk[858], n_n101, n_n1036, x128x, x5467x, x6343x}, x5482x);
	defparam lut_2936.LUT_SIZE = 6;
	defparam lut_2936.mask = 64'h00ffffffbbffbfff;

	lut_sub lut_2941 ({sk[859], i_8_, n_n38, n_n1153, x110x, x175x}, x5499x);
	defparam lut_2941.LUT_SIZE = 6;
	defparam lut_2941.mask = 64'h00ffffff0f1f0f0f;

	lut_sub lut_2944 ({sk[860], i_5_, i_2_, n_n101, x54x, x175x}, x5518x);
	defparam lut_2944.LUT_SIZE = 6;
	defparam lut_2944.mask = 64'h00ffffff00010100;

	lut_sub lut_2947 ({sk[861], i_3_, x109x, x78x, x129x, x174x}, x5519x);
	defparam lut_2947.LUT_SIZE = 6;
	defparam lut_2947.mask = 64'h00ffffff05370505;

	lut_sub lut_2950 ({sk[862], n_n58, n_n100, n_n102, n_n63, n_n77}, x5522x);
	defparam lut_2950.LUT_SIZE = 6;
	defparam lut_2950.mask = 64'h00ffffff00030057;

	lut_sub lut_2953 ({sk[863], n_n64, n_n52, x65x, x166x, x869x}, x5526x);
	defparam lut_2953.LUT_SIZE = 6;
	defparam lut_2953.mask = 64'h00ffffff7777777f;

	lut_sub lut_2957 ({sk[864], n_n78, n_n1259, x53x, n_n1176, n_n1184}, x5528x);
	defparam lut_2957.LUT_SIZE = 6;
	defparam lut_2957.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_2962 ({sk[865], n_n101, n_n100, n_n74, x340x, x5518x}, x5529x);
	defparam lut_2962.LUT_SIZE = 6;
	defparam lut_2962.mask = 64'h00ffffff7777777f;

	lut_sub lut_2966 ({sk[866], i_5_, i_3_, i_4_, x48x, x5522x}, x5531x);
	defparam lut_2966.LUT_SIZE = 6;
	defparam lut_2966.mask = 64'h00ffffff55755557;

	lut_sub lut_2970 ({sk[867], i_8_, i_6_, n_n103, n_n77, n_n1059}, x5568x);
	defparam lut_2970.LUT_SIZE = 6;
	defparam lut_2970.mask = 64'h00ffffff55555557;

	lut_sub lut_2973 ({sk[868], n_n38, n_n70, x29x, n_n1087, x153x}, x5571x);
	defparam lut_2973.LUT_SIZE = 6;
	defparam lut_2973.mask = 64'h00ffffff7777777f;

	lut_sub lut_2977 ({sk[869], n_n78, x42x, n_n1093, n_n1057, n_n1045}, x5573x);
	defparam lut_2977.LUT_SIZE = 6;
	defparam lut_2977.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2982 ({sk[870], n_n91, x53x, n_n1101, n_n1060, n_n1100}, x5574x);
	defparam lut_2982.LUT_SIZE = 6;
	defparam lut_2982.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_2987 ({sk[871], n_n77, n_n1046, x132x, n_n954, n_n939}, x5575x);
	defparam lut_2987.LUT_SIZE = 6;
	defparam lut_2987.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_2992 ({sk[872], n_n74, n_n1058, n_n971, x107x, n_n1037}, x5576x);
	defparam lut_2992.LUT_SIZE = 6;
	defparam lut_2992.mask = 64'h00ffffff5fff7fff;

	lut_sub lut_2997 ({sk[873], n_n95, x29x, x829x, x292x, n_n947}, x5579x);
	defparam lut_2997.LUT_SIZE = 6;
	defparam lut_2997.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_3002 ({sk[874], x254x, x285x, x68x, x138x}, x5580x);
	defparam lut_3002.LUT_SIZE = 5;
	defparam lut_3002.mask = 32'h0f0f7fff;

	lut_sub lut_3007 ({sk[875], x97x, x298x, x903x, x5492x, x125x}, x6358x);
	defparam lut_3007.LUT_SIZE = 6;
	defparam lut_3007.mask = 64'h00ffffff80000000;

	lut_sub lut_3009 ({sk[876], i_7_, i_8_, i_2_, x175x, x130x}, x5595x);
	defparam lut_3009.LUT_SIZE = 6;
	defparam lut_3009.mask = 64'h00ffffff01100000;

	lut_sub lut_3012 ({sk[877], n_n95, n_n1134, n_n1132, x128x, n_n962}, x5641x);
	defparam lut_3012.LUT_SIZE = 6;
	defparam lut_3012.mask = 64'h00ffffff5fff7fff;

	lut_sub lut_3017 ({sk[878], n_n101, n_n100, x78x, x128x, x218x}, x5642x);
	defparam lut_3017.LUT_SIZE = 6;
	defparam lut_3017.mask = 64'h00ffffff555f777f;

	lut_sub lut_3021 ({sk[879], n_n101, n_n1058, n_n1101, x44x, n_n954}, x5643x);
	defparam lut_3021.LUT_SIZE = 6;
	defparam lut_3021.mask = 64'h00ffffff5fff7fff;

	lut_sub lut_3026 ({sk[880], n_n1079, x324x, n_n67, x345x, n_n978}, x5644x);
	defparam lut_3026.LUT_SIZE = 6;
	defparam lut_3026.mask = 64'h00ffffff777fffff;

	lut_sub lut_3031 ({sk[881], i_1_, n_n91, x45x, n_n77, n_n959}, x6341x);
	defparam lut_3031.LUT_SIZE = 6;
	defparam lut_3031.mask = 64'h00ffffffaaa0aa80;

	lut_sub lut_3035 ({sk[882], i_7_, i_8_, n_n94, n_n66, x6341x}, x5645x);
	defparam lut_3035.LUT_SIZE = 6;
	defparam lut_3035.mask = 64'h00ffffffaaaaaaab;

	lut_sub lut_3038 ({sk[883], n_n73, n_n70, x53x, x33x, x287x}, x5646x);
	defparam lut_3038.LUT_SIZE = 6;
	defparam lut_3038.mask = 64'h00ffffff55775f7f;

	lut_sub lut_3042 ({sk[884], n_n944, n_n939, x162x, x91x, x266x}, x5648x);
	defparam lut_3042.LUT_SIZE = 6;
	defparam lut_3042.mask = 64'h00ffffff7fffffff;

	lut_sub lut_3048 ({sk[885], x1483x, x1484x, x279x, x153x, x204x}, x6340x);
	defparam lut_3048.LUT_SIZE = 6;
	defparam lut_3048.mask = 64'h00ffffff80000000;

	lut_sub lut_3050 ({sk[886], i_5_, i_3_, n_n38, n_n94, x235x}, x5664x);
	defparam lut_3050.LUT_SIZE = 6;
	defparam lut_3050.mask = 64'h00ffffff55555755;

	lut_sub lut_3053 ({sk[887], i_5_, i_3_, i_4_, n_n91, n_n94}, x5668x);
	defparam lut_3053.LUT_SIZE = 6;
	defparam lut_3053.mask = 64'h00ffffff10110000;

	lut_sub lut_3056 ({sk[888], n_n101, x55x, x112x, n_n1163, x1143x}, x5672x);
	defparam lut_3056.LUT_SIZE = 6;
	defparam lut_3056.mask = 64'h00ffffff77777fff;

	lut_sub lut_3061 ({sk[889], n_n78, x63x, x52x, n_n1216, n_n1146}, x5673x);
	defparam lut_3061.LUT_SIZE = 6;
	defparam lut_3061.mask = 64'h00ffffff77777fff;

	lut_sub lut_3066 ({sk[890], n_n94, n_n1188, n_n1193, x342x, x5493x}, x6342x);
	defparam lut_3066.LUT_SIZE = 6;
	defparam lut_3066.mask = 64'h00ffffffc0008000;

	lut_sub lut_3069 ({sk[891], i_5_, i_6_, i_3_, x328x, x350x}, x5693x);
	defparam lut_3069.LUT_SIZE = 6;
	defparam lut_3069.mask = 64'h00ffffff55557555;

	lut_sub lut_3072 ({sk[892], n_n75, n_n94, x38x, x174x, x130x}, x5694x);
	defparam lut_3072.LUT_SIZE = 6;
	defparam lut_3072.mask = 64'h00ffffff03030357;

	lut_sub lut_3075 ({sk[893], i_3_, x341x, x66x, x131x, x107x}, x5695x);
	defparam lut_3075.LUT_SIZE = 6;
	defparam lut_3075.mask = 64'h00ffffff03030357;

	lut_sub lut_3078 ({sk[894], i_5_, n_n91, x54x, x21x, x20x}, x5697x);
	defparam lut_3078.LUT_SIZE = 6;
	defparam lut_3078.mask = 64'h00ffffff05370033;

	lut_sub lut_3081 ({sk[895], i_3_, i_1_, i_2_, x333x, x339x}, x5715x);
	defparam lut_3081.LUT_SIZE = 6;
	defparam lut_3081.mask = 64'h00ffffff33333733;

	lut_sub lut_3084 ({sk[896], i_7_, i_8_, i_6_, x39x, x64x}, x6353x);
	defparam lut_3084.LUT_SIZE = 6;
	defparam lut_3084.mask = 64'h00fffffffafcffff;

	lut_sub lut_3090 ({sk[897], x255x, x226x, x71x, x876x, x877x}, x5727x);
	defparam lut_3090.LUT_SIZE = 6;
	defparam lut_3090.mask = 64'h00ffffff7fffffff;

	lut_sub lut_3096 ({sk[898], n_n1134, n_n1331, x248x, x5686x, x5687x}, x6336x);
	defparam lut_3096.LUT_SIZE = 6;
	defparam lut_3096.mask = 64'h00ffffffe0000000;

	lut_sub lut_3099 ({sk[899], i_0_, n_n91, x64x, x38x, x30x}, x5751x);
	defparam lut_3099.LUT_SIZE = 6;
	defparam lut_3099.mask = 64'h00ffffff000f111f;

	lut_sub lut_3102 ({sk[900], i_6_, i_3_, i_4_, x236x, x66x}, x5753x);
	defparam lut_3102.LUT_SIZE = 6;
	defparam lut_3102.mask = 64'h00ffffff33333373;

	lut_sub lut_3105 ({sk[901], i_7_, i_8_, x245x, x67x, n_n66}, x5758x);
	defparam lut_3105.LUT_SIZE = 6;
	defparam lut_3105.mask = 64'h00ffffff05053300;

	lut_sub lut_3108 ({sk[902], n_n91, n_n102, n_n97, n_n939, x161x}, x5763x);
	defparam lut_3108.LUT_SIZE = 6;
	defparam lut_3108.mask = 64'h00ffffff7777777f;

	lut_sub lut_3112 ({sk[903], n_n101, n_n84, n_n85, x97x, x5758x}, x5769x);
	defparam lut_3112.LUT_SIZE = 6;
	defparam lut_3112.mask = 64'h00ffffff7777777f;

	lut_sub lut_3116 ({sk[904], x256x, x215x, x141x, x142x}, x5770x);
	defparam lut_3116.LUT_SIZE = 5;
	defparam lut_3116.mask = 32'h0f0f7fff;

	lut_sub lut_3121 ({sk[905], n_n58, n_n95, n_n1132, x44x, n_n971}, x6338x);
	defparam lut_3121.LUT_SIZE = 6;
	defparam lut_3121.mask = 64'h00ffffffa0808080;

	lut_sub lut_3124 ({sk[906], x55x, n_n95, n_n983, x354x, x4944x}, x6350x);
	defparam lut_3124.LUT_SIZE = 6;
	defparam lut_3124.mask = 64'h00ffffffe0e0e000;

	lut_sub lut_3129 ({sk[907], n_n1087, x805x, x79x, x91x, x103x}, x6337x);
	defparam lut_3129.LUT_SIZE = 6;
	defparam lut_3129.mask = 64'h00ffffff80000000;

	lut_sub lut_3131 ({sk[908], i_1_, n_n80, n_n58, x110x, x234x}, x5798x);
	defparam lut_3131.LUT_SIZE = 6;
	defparam lut_3131.mask = 64'h00ffffff00550357;

	lut_sub lut_3134 ({sk[909], n_n78, x42x, n_n989, x5798x}, x5808x);
	defparam lut_3134.LUT_SIZE = 5;
	defparam lut_3134.mask = 32'h0f0f777f;

	lut_sub lut_3138 ({sk[910], x64x, n_n95, n_n969, n_n999, n_n1004}, x5809x);
	defparam lut_3138.LUT_SIZE = 6;
	defparam lut_3138.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_3143 ({sk[911], x25x, n_n95, x173x, x168x, x237x}, x5810x);
	defparam lut_3143.LUT_SIZE = 6;
	defparam lut_3143.mask = 64'h00ffffff33773f7f;

	lut_sub lut_3147 ({sk[912], n_n980, n_n983, n_n986, x753x, x5609x}, x5812x);
	defparam lut_3147.LUT_SIZE = 6;
	defparam lut_3147.mask = 64'h00ffffff7fffffff;

	lut_sub lut_3153 ({sk[913], n_n973, x145x, n_n975, x272x, x147x}, x5814x);
	defparam lut_3153.LUT_SIZE = 6;
	defparam lut_3153.mask = 64'h00ffffff7fffffff;

	lut_sub lut_3159 ({sk[914], x97x, x125x, n_n994, x163x, n_n978}, x6357x);
	defparam lut_3159.LUT_SIZE = 6;
	defparam lut_3159.mask = 64'h00ffffff80000000;

	lut_sub lut_3161 ({sk[915], n_n75, n_n74, x63x, n_n67, x5828x}, x5835x);
	defparam lut_3161.LUT_SIZE = 6;
	defparam lut_3161.mask = 64'h00ffffff00440f4f;

	lut_sub lut_3164 ({sk[916], n_n1092, n_n1091, n_n1100, x354x, x4944x}, x6335x);
	defparam lut_3164.LUT_SIZE = 6;
	defparam lut_3164.mask = 64'h00ffffffe0000000;

	lut_sub lut_3167 ({sk[917], i_5_, i_3_, i_4_, n_n78, n_n90}, x5848x);
	defparam lut_3167.LUT_SIZE = 6;
	defparam lut_3167.mask = 64'h00ffffff00100010;

	lut_sub lut_3170 ({sk[918], i_7_, i_8_, i_6_, x128x, n_n1177}, x5850x);
	defparam lut_3170.LUT_SIZE = 6;
	defparam lut_3170.mask = 64'h00ffffff55575555;

	lut_sub lut_3173 ({sk[919], i_5_, i_6_, i_3_, x316x, x344x}, x5852x);
	defparam lut_3173.LUT_SIZE = 6;
	defparam lut_3173.mask = 64'h00ffffff55555557;

	lut_sub lut_3176 ({sk[920], i_7_, i_8_, n_n103, n_n85, n_n76}, x5853x);
	defparam lut_3176.LUT_SIZE = 6;
	defparam lut_3176.mask = 64'h00ffffff05000011;

	lut_sub lut_3179 ({sk[921], i_7_, i_8_, i_6_, x239x, x41x}, x5854x);
	defparam lut_3179.LUT_SIZE = 6;
	defparam lut_3179.mask = 64'h00ffffff00530500;

	lut_sub lut_3183 ({sk[922], i_7_, i_8_, i_6_, x45x, x49x}, x5855x);
	defparam lut_3183.LUT_SIZE = 6;
	defparam lut_3183.mask = 64'h00ffffff00305000;

	lut_sub lut_3186 ({sk[923], i_5_, n_n91, n_n100, x39x, x54x}, x5856x);
	defparam lut_3186.LUT_SIZE = 6;
	defparam lut_3186.mask = 64'h00ffffff00330037;

	lut_sub lut_3189 ({sk[924], x57x, n_n92, n_n95, x88x, x132x}, x5858x);
	defparam lut_3189.LUT_SIZE = 6;
	defparam lut_3189.mask = 64'h00ffffff33773f7f;

	lut_sub lut_3193 ({sk[925], i_5_, x54x, x343x, x48x, x185x}, x5859x);
	defparam lut_3193.LUT_SIZE = 6;
	defparam lut_3193.mask = 64'h00ffffff5f5f5f7f;

	lut_sub lut_3197 ({sk[926], n_n73, x111x, n_n1169, x120x, x238x}, x5860x);
	defparam lut_3197.LUT_SIZE = 6;
	defparam lut_3197.mask = 64'h00ffffff3f3f3f7f;

	lut_sub lut_3201 ({sk[927], n_n52, n_n82, x21x, x22x, x5856x}, x5866x);
	defparam lut_3201.LUT_SIZE = 6;
	defparam lut_3201.mask = 64'h00ffffff555f777f;

	lut_sub lut_3205 ({sk[928], i_2_, x55x, n_n95, x5493x, x175x}, x5880x);
	defparam lut_3205.LUT_SIZE = 6;
	defparam lut_3205.mask = 64'h00ffffff111f000f;

	lut_sub lut_3208 ({sk[929], i_7_, i_8_, i_3_, x5687x, n_n1009}, x5881x);
	defparam lut_3208.LUT_SIZE = 6;
	defparam lut_3208.mask = 64'h00ffffff75555555;

	lut_sub lut_3211 ({sk[930], i_3_, i_1_, i_2_, x339x, n_n1013}, x5882x);
	defparam lut_3211.LUT_SIZE = 6;
	defparam lut_3211.mask = 64'h00ffffff55555755;

	lut_sub lut_3214 ({sk[931], n_n81, n_n91, n_n103, n_n102, n_n82}, x5899x);
	defparam lut_3214.LUT_SIZE = 6;
	defparam lut_3214.mask = 64'h00ffffff00030507;

	lut_sub lut_3217 ({sk[932], i_3_, i_1_, i_2_, x78x, x324x}, x5914x);
	defparam lut_3217.LUT_SIZE = 6;
	defparam lut_3217.mask = 64'h00ffffff00050300;

	lut_sub lut_3220 ({sk[933], n_n93, n_n103, n_n74, x38x, x174x}, x5915x);
	defparam lut_3220.LUT_SIZE = 6;
	defparam lut_3220.mask = 64'h00ffffff1111111f;

	lut_sub lut_3223 ({sk[934], i_3_, n_n58, x19x, x109x, x20x}, x5918x);
	defparam lut_3223.LUT_SIZE = 6;
	defparam lut_3223.mask = 64'h00ffffff000f111f;

	lut_sub lut_3226 ({sk[935], i_5_, x32x, x54x, x346x, x190x}, x5919x);
	defparam lut_3226.LUT_SIZE = 6;
	defparam lut_3226.mask = 64'h00ffffff7777777f;

	lut_sub lut_3230 ({sk[936], n_n58, x26x, x32x, n_n102, x157x}, x5921x);
	defparam lut_3230.LUT_SIZE = 6;
	defparam lut_3230.mask = 64'h00ffffff575757ff;

	lut_sub lut_3234 ({sk[937], n_n78, n_n92, n_n85, x210x, x663x}, x5922x);
	defparam lut_3234.LUT_SIZE = 6;
	defparam lut_3234.mask = 64'h00ffffff7777777f;

	lut_sub lut_3238 ({sk[938], x235x, n_n1286, x131x, x5068x, n_n1158}, x5924x);
	defparam lut_3238.LUT_SIZE = 6;
	defparam lut_3238.mask = 64'h00ffffff57ffffff;

	lut_sub lut_3243 ({sk[939], n_n75, x45x, x25x, n_n95, x5915x}, x5926x);
	defparam lut_3243.LUT_SIZE = 6;
	defparam lut_3243.mask = 64'h00ffffff55775f7f;

	lut_sub lut_3247 ({sk[940], n_n52, n_n101, x21x, x22x, x5918x}, x5927x);
	defparam lut_3247.LUT_SIZE = 6;
	defparam lut_3247.mask = 64'h00ffffff555f777f;

	lut_sub lut_3251 ({sk[941], n_n1312, x129x, x5338x, x5914x, x5926x}, x5933x);
	defparam lut_3251.LUT_SIZE = 6;
	defparam lut_3251.mask = 64'h00ffffff777fffff;

	lut_sub lut_3256 ({sk[942], i_5_, i_4_, n_n58, n_n1039, x327x}, x5944x);
	defparam lut_3256.LUT_SIZE = 6;
	defparam lut_3256.mask = 64'h00ffffff37333333;

	lut_sub lut_3259 ({sk[943], i_6_, i_3_, i_4_, x66x, n_n1013}, x5946x);
	defparam lut_3259.LUT_SIZE = 6;
	defparam lut_3259.mask = 64'h00ffffff55555575;

	lut_sub lut_3262 ({sk[944], i_5_, n_n80, x337x, x247x, x28x}, x5965x);
	defparam lut_3262.LUT_SIZE = 6;
	defparam lut_3262.mask = 64'h00ffffff111f000f;

	lut_sub lut_3265 ({sk[945], n_n64, n_n100, x25x, n_n76, x247x}, x5966x);
	defparam lut_3265.LUT_SIZE = 6;
	defparam lut_3265.mask = 64'h00ffffff05050537;

	lut_sub lut_3268 ({sk[946], i_3_, x19x, x109x, x177x, x129x}, x5967x);
	defparam lut_3268.LUT_SIZE = 6;
	defparam lut_3268.mask = 64'h00ffffff05370033;

	lut_sub lut_3271 ({sk[947], i_6_, x76x, n_n63, x110x, x66x}, x5968x);
	defparam lut_3271.LUT_SIZE = 6;
	defparam lut_3271.mask = 64'h00ffffff000f111f;

	lut_sub lut_3274 ({sk[948], n_n101, n_n100, n_n102, n_n63, n_n90}, x5969x);
	defparam lut_3274.LUT_SIZE = 6;
	defparam lut_3274.mask = 64'h00ffffff0101010f;

	lut_sub lut_3277 ({sk[949], i_5_, i_3_, i_4_, x88x, x20x}, x5971x);
	defparam lut_3277.LUT_SIZE = 6;
	defparam lut_3277.mask = 64'h00ffffff33333337;

	lut_sub lut_3280 ({sk[950], n_n78, x27x, n_n1193, x1291x, x1292x}, x5972x);
	defparam lut_3280.LUT_SIZE = 6;
	defparam lut_3280.mask = 64'h00ffffff7f7f7fff;

	lut_sub lut_3285 ({sk[951], n_n78, n_n102, n_n85, n_n1297, x220x}, x5974x);
	defparam lut_3285.LUT_SIZE = 6;
	defparam lut_3285.mask = 64'h00ffffff7777777f;

	lut_sub lut_3289 ({sk[952], n_n81, n_n92, x32x, x37x, x5969x}, x6360x);
	defparam lut_3289.LUT_SIZE = 6;
	defparam lut_3289.mask = 64'h00ffffffaaa08080;

	lut_sub lut_3293 ({sk[953], i_8_, i_4_, n_n38, n_n1092, x242x}, x5996x);
	defparam lut_3293.LUT_SIZE = 6;
	defparam lut_3293.mask = 64'h00ffffff37333333;

	lut_sub lut_3296 ({sk[954], i_2_, n_n101, n_n78, n_n77, x108x}, x6006x);
	defparam lut_3296.LUT_SIZE = 6;
	defparam lut_3296.mask = 64'h00ffffff00110303;

	lut_sub lut_3299 ({sk[955], n_n91, n_n102, n_n97, n_n939, x268x}, x6009x);
	defparam lut_3299.LUT_SIZE = 6;
	defparam lut_3299.mask = 64'h00ffffff7777777f;

	lut_sub lut_3303 ({sk[956], n_n101, n_n74, n_n90, x94x, x1348x}, x6010x);
	defparam lut_3303.LUT_SIZE = 6;
	defparam lut_3303.mask = 64'h00ffffff7777777f;

	lut_sub lut_3307 ({sk[957], n_n86, n_n97, n_n77, n_n1128, x5996x}, x6011x);
	defparam lut_3307.LUT_SIZE = 6;
	defparam lut_3307.mask = 64'h00ffffff7777777f;

	lut_sub lut_3311 ({sk[958], n_n83, x251x, x321x, n_n1176, x320x}, x6012x);
	defparam lut_3311.LUT_SIZE = 6;
	defparam lut_3311.mask = 64'h00ffffff3fff7fff;

	lut_sub lut_3316 ({sk[959], n_n969, n_n1184, n_n1156, x5686x, x5687x}, x6013x);
	defparam lut_3316.LUT_SIZE = 6;
	defparam lut_3316.mask = 64'h00ffffff1fffffff;

	lut_sub lut_3321 ({sk[960], n_n78, n_n941, x237x, n_n1164, n_n975}, x6014x);
	defparam lut_3321.LUT_SIZE = 6;
	defparam lut_3321.mask = 64'h00ffffff77ff7fff;

	lut_sub lut_3326 ({sk[961], n_n91, x63x, x83x, x22x, n_n966}, x6015x);
	defparam lut_3326.LUT_SIZE = 6;
	defparam lut_3326.mask = 64'h00ffffff55557fff;

	lut_sub lut_3331 ({sk[962], i_7_, i_6_, x21x, x336x, x6006x}, x6016x);
	defparam lut_3331.LUT_SIZE = 6;
	defparam lut_3331.mask = 64'h00ffffff777f7777;

	lut_sub lut_3335 ({sk[963], n_n70, x53x, x215x, x150x, x153x}, x6018x);
	defparam lut_3335.LUT_SIZE = 6;
	defparam lut_3335.mask = 64'h00ffffff7f7f7fff;


endmodule